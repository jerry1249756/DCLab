
module Altpll (
	reset_reset_n,
	clk_clk,
	altpll_0_c0_clk,
	altpll_1_c0_clk);	

	input		reset_reset_n;
	input		clk_clk;
	output		altpll_0_c0_clk;
	output		altpll_1_c0_clk;
endmodule
