
module Altpll (
	altpll_0_c25m_clk,
	altpll_0_c3p2m_clk,
	altpll_0_c50k_clk,
	clk_clk,
	reset_reset_n);	

	output		altpll_0_c25m_clk;
	output		altpll_0_c3p2m_clk;
	output		altpll_0_c50k_clk;
	input		clk_clk;
	input		reset_reset_n;
endmodule
