module Coordinate_generator(
    input signed [$clog2(`PIXEL_COLUMN)-1:0] p_x,  //-39~39
    input signed [$clog2(`PIXEL_ROW)-1:0] p_y,     //-29~29
    output signed [6:0] real_x[15:0],
    output signed [6:0] real_y[15:0]
);
    logic signed [$clog2(`PIXEL_COLUMN)-1:0] temp_x;
    logic signed [$clog2(`PIXEL_ROW)-1:0] temp_y;
    assign temp_x = (p_x==-40) ? p_x+1 : p_x;
    assign temp_y = (p_y==-30) ? p_y+1 : p_y;
    genvar idx;
    generate
        for(idx=0; idx<4; idx=idx+1) begin: Geny1
            assign real_y[idx] = temp_y + 15;
        end
        for(idx=4; idx<8; idx=idx+1) begin: Geny2
            assign real_y[idx] = temp_y + 5;
        end
        for(idx=8; idx<12; idx=idx+1) begin: Geny3
            assign real_y[idx] = temp_y - 5;
        end
        for(idx=12; idx<16; idx=idx+1) begin: Geny4
            assign real_y[idx] = temp_y - 15;
        end
        for(idx=0; idx<16; idx=idx+4) begin: Genx1
            assign real_x[idx] = temp_x + 15;
        end
        for(idx=1; idx<16; idx=idx+4) begin: Genx2
            assign real_x[idx] = temp_x + 5;
        end
        for(idx=2; idx<16; idx=idx+4) begin:Genx3
            assign real_x[idx] = temp_x - 5;
        end
        for(idx=3; idx<16; idx=idx+4) begin:Genx4
            assign real_x[idx] = temp_x - 15;
        end
    endgenerate
endmodule

module abs_X(
    input signed [6:0] x,
    output [6:0] abs_real_x
);
    assign abs_real_x = x[6] ? -x : x;
endmodule

module abs_Y(
    input signed [6:0] y,
    output [6:0] abs_real_y
);
    assign abs_real_y = y[6] ? -y : y;
endmodule

module Delta_generator (
    input signed [$clog2(`PIXEL_COLUMN)-1:0] p_x,
    input signed [$clog2(`PIXEL_ROW)-1:0] p_y,
    output [6:0] delta[15:0]
);
    logic signed [6:0] real_x[15:0];
    logic signed [6:0] real_y[15:0];
    logic [6:0] abs_real_x[15:0];
    logic [6:0] abs_real_y[15:0];
    logic [5:0] data [2474:0];

    assign data[0] = 6'b000000;
    assign data[1] = 6'b000000;
    assign data[2] = 6'b000000;
    assign data[3] = 6'b000000;
    assign data[4] = 6'b000000;
    assign data[5] = 6'b000000;
    assign data[6] = 6'b000000;
    assign data[7] = 6'b000000;
    assign data[8] = 6'b000001;
    assign data[9] = 6'b000001;
    assign data[10] = 6'b000001;
    assign data[11] = 6'b000001;
    assign data[12] = 6'b000010;
    assign data[13] = 6'b000010;
    assign data[14] = 6'b000011;
    assign data[15] = 6'b000011;
    assign data[16] = 6'b000011;
    assign data[17] = 6'b000100;
    assign data[18] = 6'b000100;
    assign data[19] = 6'b000101;
    assign data[20] = 6'b000101;
    assign data[21] = 6'b000110;
    assign data[22] = 6'b000111;
    assign data[23] = 6'b000111;
    assign data[24] = 6'b001000;
    assign data[25] = 6'b001001;
    assign data[26] = 6'b001001;
    assign data[27] = 6'b001010;
    assign data[28] = 6'b001011;
    assign data[29] = 6'b001011;
    assign data[30] = 6'b001100;
    assign data[31] = 6'b001101;
    assign data[32] = 6'b001110;
    assign data[33] = 6'b001111;
    assign data[34] = 6'b001111;
    assign data[35] = 6'b010000;
    assign data[36] = 6'b010001;
    assign data[37] = 6'b010010;
    assign data[38] = 6'b010011;
    assign data[39] = 6'b010100;
    assign data[40] = 6'b010101;
    assign data[41] = 6'b010110;
    assign data[42] = 6'b010111;
    assign data[43] = 6'b010111;
    assign data[44] = 6'b011000;
    assign data[45] = 6'b000000;
    assign data[46] = 6'b000000;
    assign data[47] = 6'b000000;
    assign data[48] = 6'b000000;
    assign data[49] = 6'b000000;
    assign data[50] = 6'b000000;
    assign data[51] = 6'b000000;
    assign data[52] = 6'b000000;
    assign data[53] = 6'b000001;
    assign data[54] = 6'b000001;
    assign data[55] = 6'b000001;
    assign data[56] = 6'b000001;
    assign data[57] = 6'b000010;
    assign data[58] = 6'b000010;
    assign data[59] = 6'b000011;
    assign data[60] = 6'b000011;
    assign data[61] = 6'b000011;
    assign data[62] = 6'b000100;
    assign data[63] = 6'b000100;
    assign data[64] = 6'b000101;
    assign data[65] = 6'b000110;
    assign data[66] = 6'b000110;
    assign data[67] = 6'b000111;
    assign data[68] = 6'b000111;
    assign data[69] = 6'b001000;
    assign data[70] = 6'b001001;
    assign data[71] = 6'b001001;
    assign data[72] = 6'b001010;
    assign data[73] = 6'b001011;
    assign data[74] = 6'b001011;
    assign data[75] = 6'b001100;
    assign data[76] = 6'b001101;
    assign data[77] = 6'b001110;
    assign data[78] = 6'b001111;
    assign data[79] = 6'b001111;
    assign data[80] = 6'b010000;
    assign data[81] = 6'b010001;
    assign data[82] = 6'b010010;
    assign data[83] = 6'b010011;
    assign data[84] = 6'b010100;
    assign data[85] = 6'b010101;
    assign data[86] = 6'b010110;
    assign data[87] = 6'b010111;
    assign data[88] = 6'b010111;
    assign data[89] = 6'b011000;
    assign data[90] = 6'b000000;
    assign data[91] = 6'b000000;
    assign data[92] = 6'b000000;
    assign data[93] = 6'b000000;
    assign data[94] = 6'b000000;
    assign data[95] = 6'b000000;
    assign data[96] = 6'b000000;
    assign data[97] = 6'b000000;
    assign data[98] = 6'b000001;
    assign data[99] = 6'b000001;
    assign data[100] = 6'b000001;
    assign data[101] = 6'b000010;
    assign data[102] = 6'b000010;
    assign data[103] = 6'b000010;
    assign data[104] = 6'b000011;
    assign data[105] = 6'b000011;
    assign data[106] = 6'b000100;
    assign data[107] = 6'b000100;
    assign data[108] = 6'b000100;
    assign data[109] = 6'b000101;
    assign data[110] = 6'b000110;
    assign data[111] = 6'b000110;
    assign data[112] = 6'b000111;
    assign data[113] = 6'b000111;
    assign data[114] = 6'b001000;
    assign data[115] = 6'b001001;
    assign data[116] = 6'b001001;
    assign data[117] = 6'b001010;
    assign data[118] = 6'b001011;
    assign data[119] = 6'b001011;
    assign data[120] = 6'b001100;
    assign data[121] = 6'b001101;
    assign data[122] = 6'b001110;
    assign data[123] = 6'b001111;
    assign data[124] = 6'b001111;
    assign data[125] = 6'b010000;
    assign data[126] = 6'b010001;
    assign data[127] = 6'b010010;
    assign data[128] = 6'b010011;
    assign data[129] = 6'b010100;
    assign data[130] = 6'b010101;
    assign data[131] = 6'b010110;
    assign data[132] = 6'b010111;
    assign data[133] = 6'b011000;
    assign data[134] = 6'b011001;
    assign data[135] = 6'b000000;
    assign data[136] = 6'b000000;
    assign data[137] = 6'b000000;
    assign data[138] = 6'b000000;
    assign data[139] = 6'b000000;
    assign data[140] = 6'b000000;
    assign data[141] = 6'b000000;
    assign data[142] = 6'b000001;
    assign data[143] = 6'b000001;
    assign data[144] = 6'b000001;
    assign data[145] = 6'b000001;
    assign data[146] = 6'b000010;
    assign data[147] = 6'b000010;
    assign data[148] = 6'b000010;
    assign data[149] = 6'b000011;
    assign data[150] = 6'b000011;
    assign data[151] = 6'b000100;
    assign data[152] = 6'b000100;
    assign data[153] = 6'b000101;
    assign data[154] = 6'b000101;
    assign data[155] = 6'b000110;
    assign data[156] = 6'b000110;
    assign data[157] = 6'b000111;
    assign data[158] = 6'b000111;
    assign data[159] = 6'b001000;
    assign data[160] = 6'b001001;
    assign data[161] = 6'b001001;
    assign data[162] = 6'b001010;
    assign data[163] = 6'b001011;
    assign data[164] = 6'b001100;
    assign data[165] = 6'b001100;
    assign data[166] = 6'b001101;
    assign data[167] = 6'b001110;
    assign data[168] = 6'b001111;
    assign data[169] = 6'b001111;
    assign data[170] = 6'b010000;
    assign data[171] = 6'b010001;
    assign data[172] = 6'b010010;
    assign data[173] = 6'b010011;
    assign data[174] = 6'b010100;
    assign data[175] = 6'b010101;
    assign data[176] = 6'b010110;
    assign data[177] = 6'b010111;
    assign data[178] = 6'b011000;
    assign data[179] = 6'b011001;
    assign data[180] = 6'b000000;
    assign data[181] = 6'b000000;
    assign data[182] = 6'b000000;
    assign data[183] = 6'b000000;
    assign data[184] = 6'b000000;
    assign data[185] = 6'b000000;
    assign data[186] = 6'b000000;
    assign data[187] = 6'b000001;
    assign data[188] = 6'b000001;
    assign data[189] = 6'b000001;
    assign data[190] = 6'b000001;
    assign data[191] = 6'b000010;
    assign data[192] = 6'b000010;
    assign data[193] = 6'b000010;
    assign data[194] = 6'b000011;
    assign data[195] = 6'b000011;
    assign data[196] = 6'b000100;
    assign data[197] = 6'b000100;
    assign data[198] = 6'b000101;
    assign data[199] = 6'b000101;
    assign data[200] = 6'b000110;
    assign data[201] = 6'b000110;
    assign data[202] = 6'b000111;
    assign data[203] = 6'b001000;
    assign data[204] = 6'b001000;
    assign data[205] = 6'b001001;
    assign data[206] = 6'b001001;
    assign data[207] = 6'b001010;
    assign data[208] = 6'b001011;
    assign data[209] = 6'b001100;
    assign data[210] = 6'b001100;
    assign data[211] = 6'b001101;
    assign data[212] = 6'b001110;
    assign data[213] = 6'b001111;
    assign data[214] = 6'b010000;
    assign data[215] = 6'b010000;
    assign data[216] = 6'b010001;
    assign data[217] = 6'b010010;
    assign data[218] = 6'b010011;
    assign data[219] = 6'b010100;
    assign data[220] = 6'b010101;
    assign data[221] = 6'b010110;
    assign data[222] = 6'b010111;
    assign data[223] = 6'b011000;
    assign data[224] = 6'b011001;
    assign data[225] = 6'b000000;
    assign data[226] = 6'b000000;
    assign data[227] = 6'b000000;
    assign data[228] = 6'b000000;
    assign data[229] = 6'b000000;
    assign data[230] = 6'b000000;
    assign data[231] = 6'b000001;
    assign data[232] = 6'b000001;
    assign data[233] = 6'b000001;
    assign data[234] = 6'b000001;
    assign data[235] = 6'b000010;
    assign data[236] = 6'b000010;
    assign data[237] = 6'b000010;
    assign data[238] = 6'b000011;
    assign data[239] = 6'b000011;
    assign data[240] = 6'b000011;
    assign data[241] = 6'b000100;
    assign data[242] = 6'b000100;
    assign data[243] = 6'b000101;
    assign data[244] = 6'b000101;
    assign data[245] = 6'b000110;
    assign data[246] = 6'b000110;
    assign data[247] = 6'b000111;
    assign data[248] = 6'b001000;
    assign data[249] = 6'b001000;
    assign data[250] = 6'b001001;
    assign data[251] = 6'b001010;
    assign data[252] = 6'b001010;
    assign data[253] = 6'b001011;
    assign data[254] = 6'b001100;
    assign data[255] = 6'b001101;
    assign data[256] = 6'b001101;
    assign data[257] = 6'b001110;
    assign data[258] = 6'b001111;
    assign data[259] = 6'b010000;
    assign data[260] = 6'b010001;
    assign data[261] = 6'b010001;
    assign data[262] = 6'b010010;
    assign data[263] = 6'b010011;
    assign data[264] = 6'b010100;
    assign data[265] = 6'b010101;
    assign data[266] = 6'b010110;
    assign data[267] = 6'b010111;
    assign data[268] = 6'b011000;
    assign data[269] = 6'b011001;
    assign data[270] = 6'b000000;
    assign data[271] = 6'b000000;
    assign data[272] = 6'b000000;
    assign data[273] = 6'b000000;
    assign data[274] = 6'b000000;
    assign data[275] = 6'b000001;
    assign data[276] = 6'b000001;
    assign data[277] = 6'b000001;
    assign data[278] = 6'b000001;
    assign data[279] = 6'b000001;
    assign data[280] = 6'b000010;
    assign data[281] = 6'b000010;
    assign data[282] = 6'b000010;
    assign data[283] = 6'b000011;
    assign data[284] = 6'b000011;
    assign data[285] = 6'b000100;
    assign data[286] = 6'b000100;
    assign data[287] = 6'b000100;
    assign data[288] = 6'b000101;
    assign data[289] = 6'b000110;
    assign data[290] = 6'b000110;
    assign data[291] = 6'b000111;
    assign data[292] = 6'b000111;
    assign data[293] = 6'b001000;
    assign data[294] = 6'b001000;
    assign data[295] = 6'b001001;
    assign data[296] = 6'b001010;
    assign data[297] = 6'b001010;
    assign data[298] = 6'b001011;
    assign data[299] = 6'b001100;
    assign data[300] = 6'b001101;
    assign data[301] = 6'b001101;
    assign data[302] = 6'b001110;
    assign data[303] = 6'b001111;
    assign data[304] = 6'b010000;
    assign data[305] = 6'b010001;
    assign data[306] = 6'b010010;
    assign data[307] = 6'b010010;
    assign data[308] = 6'b010011;
    assign data[309] = 6'b010100;
    assign data[310] = 6'b010101;
    assign data[311] = 6'b010110;
    assign data[312] = 6'b010111;
    assign data[313] = 6'b011000;
    assign data[314] = 6'b011001;
    assign data[315] = 6'b000000;
    assign data[316] = 6'b000000;
    assign data[317] = 6'b000000;
    assign data[318] = 6'b000001;
    assign data[319] = 6'b000001;
    assign data[320] = 6'b000001;
    assign data[321] = 6'b000001;
    assign data[322] = 6'b000001;
    assign data[323] = 6'b000001;
    assign data[324] = 6'b000010;
    assign data[325] = 6'b000010;
    assign data[326] = 6'b000010;
    assign data[327] = 6'b000011;
    assign data[328] = 6'b000011;
    assign data[329] = 6'b000011;
    assign data[330] = 6'b000100;
    assign data[331] = 6'b000100;
    assign data[332] = 6'b000101;
    assign data[333] = 6'b000101;
    assign data[334] = 6'b000110;
    assign data[335] = 6'b000110;
    assign data[336] = 6'b000111;
    assign data[337] = 6'b000111;
    assign data[338] = 6'b001000;
    assign data[339] = 6'b001001;
    assign data[340] = 6'b001001;
    assign data[341] = 6'b001010;
    assign data[342] = 6'b001011;
    assign data[343] = 6'b001011;
    assign data[344] = 6'b001100;
    assign data[345] = 6'b001101;
    assign data[346] = 6'b001110;
    assign data[347] = 6'b001110;
    assign data[348] = 6'b001111;
    assign data[349] = 6'b010000;
    assign data[350] = 6'b010001;
    assign data[351] = 6'b010010;
    assign data[352] = 6'b010011;
    assign data[353] = 6'b010011;
    assign data[354] = 6'b010100;
    assign data[355] = 6'b010101;
    assign data[356] = 6'b010110;
    assign data[357] = 6'b010111;
    assign data[358] = 6'b011000;
    assign data[359] = 6'b011001;
    assign data[360] = 6'b000001;
    assign data[361] = 6'b000001;
    assign data[362] = 6'b000001;
    assign data[363] = 6'b000001;
    assign data[364] = 6'b000001;
    assign data[365] = 6'b000001;
    assign data[366] = 6'b000001;
    assign data[367] = 6'b000001;
    assign data[368] = 6'b000010;
    assign data[369] = 6'b000010;
    assign data[370] = 6'b000010;
    assign data[371] = 6'b000010;
    assign data[372] = 6'b000011;
    assign data[373] = 6'b000011;
    assign data[374] = 6'b000100;
    assign data[375] = 6'b000100;
    assign data[376] = 6'b000100;
    assign data[377] = 6'b000101;
    assign data[378] = 6'b000101;
    assign data[379] = 6'b000110;
    assign data[380] = 6'b000110;
    assign data[381] = 6'b000111;
    assign data[382] = 6'b001000;
    assign data[383] = 6'b001000;
    assign data[384] = 6'b001001;
    assign data[385] = 6'b001001;
    assign data[386] = 6'b001010;
    assign data[387] = 6'b001011;
    assign data[388] = 6'b001100;
    assign data[389] = 6'b001100;
    assign data[390] = 6'b001101;
    assign data[391] = 6'b001110;
    assign data[392] = 6'b001111;
    assign data[393] = 6'b001111;
    assign data[394] = 6'b010000;
    assign data[395] = 6'b010001;
    assign data[396] = 6'b010010;
    assign data[397] = 6'b010011;
    assign data[398] = 6'b010100;
    assign data[399] = 6'b010101;
    assign data[400] = 6'b010101;
    assign data[401] = 6'b010110;
    assign data[402] = 6'b010111;
    assign data[403] = 6'b011000;
    assign data[404] = 6'b011001;
    assign data[405] = 6'b000001;
    assign data[406] = 6'b000001;
    assign data[407] = 6'b000001;
    assign data[408] = 6'b000001;
    assign data[409] = 6'b000001;
    assign data[410] = 6'b000001;
    assign data[411] = 6'b000001;
    assign data[412] = 6'b000010;
    assign data[413] = 6'b000010;
    assign data[414] = 6'b000010;
    assign data[415] = 6'b000010;
    assign data[416] = 6'b000011;
    assign data[417] = 6'b000011;
    assign data[418] = 6'b000011;
    assign data[419] = 6'b000100;
    assign data[420] = 6'b000100;
    assign data[421] = 6'b000101;
    assign data[422] = 6'b000101;
    assign data[423] = 6'b000110;
    assign data[424] = 6'b000110;
    assign data[425] = 6'b000111;
    assign data[426] = 6'b000111;
    assign data[427] = 6'b001000;
    assign data[428] = 6'b001000;
    assign data[429] = 6'b001001;
    assign data[430] = 6'b001010;
    assign data[431] = 6'b001010;
    assign data[432] = 6'b001011;
    assign data[433] = 6'b001100;
    assign data[434] = 6'b001101;
    assign data[435] = 6'b001101;
    assign data[436] = 6'b001110;
    assign data[437] = 6'b001111;
    assign data[438] = 6'b010000;
    assign data[439] = 6'b010000;
    assign data[440] = 6'b010001;
    assign data[441] = 6'b010010;
    assign data[442] = 6'b010011;
    assign data[443] = 6'b010100;
    assign data[444] = 6'b010101;
    assign data[445] = 6'b010110;
    assign data[446] = 6'b010111;
    assign data[447] = 6'b011000;
    assign data[448] = 6'b011000;
    assign data[449] = 6'b011001;
    assign data[450] = 6'b000001;
    assign data[451] = 6'b000001;
    assign data[452] = 6'b000001;
    assign data[453] = 6'b000001;
    assign data[454] = 6'b000001;
    assign data[455] = 6'b000010;
    assign data[456] = 6'b000010;
    assign data[457] = 6'b000010;
    assign data[458] = 6'b000010;
    assign data[459] = 6'b000010;
    assign data[460] = 6'b000011;
    assign data[461] = 6'b000011;
    assign data[462] = 6'b000011;
    assign data[463] = 6'b000100;
    assign data[464] = 6'b000100;
    assign data[465] = 6'b000101;
    assign data[466] = 6'b000101;
    assign data[467] = 6'b000101;
    assign data[468] = 6'b000110;
    assign data[469] = 6'b000110;
    assign data[470] = 6'b000111;
    assign data[471] = 6'b001000;
    assign data[472] = 6'b001000;
    assign data[473] = 6'b001001;
    assign data[474] = 6'b001001;
    assign data[475] = 6'b001010;
    assign data[476] = 6'b001011;
    assign data[477] = 6'b001011;
    assign data[478] = 6'b001100;
    assign data[479] = 6'b001101;
    assign data[480] = 6'b001110;
    assign data[481] = 6'b001110;
    assign data[482] = 6'b001111;
    assign data[483] = 6'b010000;
    assign data[484] = 6'b010001;
    assign data[485] = 6'b010001;
    assign data[486] = 6'b010010;
    assign data[487] = 6'b010011;
    assign data[488] = 6'b010100;
    assign data[489] = 6'b010101;
    assign data[490] = 6'b010110;
    assign data[491] = 6'b010111;
    assign data[492] = 6'b011000;
    assign data[493] = 6'b011001;
    assign data[494] = 6'b011010;
    assign data[495] = 6'b000001;
    assign data[496] = 6'b000001;
    assign data[497] = 6'b000010;
    assign data[498] = 6'b000010;
    assign data[499] = 6'b000010;
    assign data[500] = 6'b000010;
    assign data[501] = 6'b000010;
    assign data[502] = 6'b000010;
    assign data[503] = 6'b000010;
    assign data[504] = 6'b000011;
    assign data[505] = 6'b000011;
    assign data[506] = 6'b000011;
    assign data[507] = 6'b000100;
    assign data[508] = 6'b000100;
    assign data[509] = 6'b000100;
    assign data[510] = 6'b000101;
    assign data[511] = 6'b000101;
    assign data[512] = 6'b000110;
    assign data[513] = 6'b000110;
    assign data[514] = 6'b000111;
    assign data[515] = 6'b000111;
    assign data[516] = 6'b001000;
    assign data[517] = 6'b001000;
    assign data[518] = 6'b001001;
    assign data[519] = 6'b001010;
    assign data[520] = 6'b001010;
    assign data[521] = 6'b001011;
    assign data[522] = 6'b001100;
    assign data[523] = 6'b001100;
    assign data[524] = 6'b001101;
    assign data[525] = 6'b001110;
    assign data[526] = 6'b001111;
    assign data[527] = 6'b001111;
    assign data[528] = 6'b010000;
    assign data[529] = 6'b010001;
    assign data[530] = 6'b010010;
    assign data[531] = 6'b010011;
    assign data[532] = 6'b010011;
    assign data[533] = 6'b010100;
    assign data[534] = 6'b010101;
    assign data[535] = 6'b010110;
    assign data[536] = 6'b010111;
    assign data[537] = 6'b011000;
    assign data[538] = 6'b011001;
    assign data[539] = 6'b011010;
    assign data[540] = 6'b000010;
    assign data[541] = 6'b000010;
    assign data[542] = 6'b000010;
    assign data[543] = 6'b000010;
    assign data[544] = 6'b000010;
    assign data[545] = 6'b000010;
    assign data[546] = 6'b000010;
    assign data[547] = 6'b000011;
    assign data[548] = 6'b000011;
    assign data[549] = 6'b000011;
    assign data[550] = 6'b000011;
    assign data[551] = 6'b000100;
    assign data[552] = 6'b000100;
    assign data[553] = 6'b000100;
    assign data[554] = 6'b000101;
    assign data[555] = 6'b000101;
    assign data[556] = 6'b000110;
    assign data[557] = 6'b000110;
    assign data[558] = 6'b000111;
    assign data[559] = 6'b000111;
    assign data[560] = 6'b001000;
    assign data[561] = 6'b001000;
    assign data[562] = 6'b001001;
    assign data[563] = 6'b001001;
    assign data[564] = 6'b001010;
    assign data[565] = 6'b001011;
    assign data[566] = 6'b001011;
    assign data[567] = 6'b001100;
    assign data[568] = 6'b001101;
    assign data[569] = 6'b001101;
    assign data[570] = 6'b001110;
    assign data[571] = 6'b001111;
    assign data[572] = 6'b010000;
    assign data[573] = 6'b010000;
    assign data[574] = 6'b010001;
    assign data[575] = 6'b010010;
    assign data[576] = 6'b010011;
    assign data[577] = 6'b010100;
    assign data[578] = 6'b010101;
    assign data[579] = 6'b010101;
    assign data[580] = 6'b010110;
    assign data[581] = 6'b010111;
    assign data[582] = 6'b011000;
    assign data[583] = 6'b011001;
    assign data[584] = 6'b011010;
    assign data[585] = 6'b000010;
    assign data[586] = 6'b000010;
    assign data[587] = 6'b000010;
    assign data[588] = 6'b000010;
    assign data[589] = 6'b000010;
    assign data[590] = 6'b000011;
    assign data[591] = 6'b000011;
    assign data[592] = 6'b000011;
    assign data[593] = 6'b000011;
    assign data[594] = 6'b000011;
    assign data[595] = 6'b000100;
    assign data[596] = 6'b000100;
    assign data[597] = 6'b000100;
    assign data[598] = 6'b000101;
    assign data[599] = 6'b000101;
    assign data[600] = 6'b000110;
    assign data[601] = 6'b000110;
    assign data[602] = 6'b000110;
    assign data[603] = 6'b000111;
    assign data[604] = 6'b000111;
    assign data[605] = 6'b001000;
    assign data[606] = 6'b001000;
    assign data[607] = 6'b001001;
    assign data[608] = 6'b001010;
    assign data[609] = 6'b001010;
    assign data[610] = 6'b001011;
    assign data[611] = 6'b001100;
    assign data[612] = 6'b001100;
    assign data[613] = 6'b001101;
    assign data[614] = 6'b001110;
    assign data[615] = 6'b001110;
    assign data[616] = 6'b001111;
    assign data[617] = 6'b010000;
    assign data[618] = 6'b010001;
    assign data[619] = 6'b010010;
    assign data[620] = 6'b010010;
    assign data[621] = 6'b010011;
    assign data[622] = 6'b010100;
    assign data[623] = 6'b010101;
    assign data[624] = 6'b010110;
    assign data[625] = 6'b010111;
    assign data[626] = 6'b011000;
    assign data[627] = 6'b011001;
    assign data[628] = 6'b011001;
    assign data[629] = 6'b011010;
    assign data[630] = 6'b000011;
    assign data[631] = 6'b000011;
    assign data[632] = 6'b000011;
    assign data[633] = 6'b000011;
    assign data[634] = 6'b000011;
    assign data[635] = 6'b000011;
    assign data[636] = 6'b000011;
    assign data[637] = 6'b000011;
    assign data[638] = 6'b000100;
    assign data[639] = 6'b000100;
    assign data[640] = 6'b000100;
    assign data[641] = 6'b000100;
    assign data[642] = 6'b000101;
    assign data[643] = 6'b000101;
    assign data[644] = 6'b000101;
    assign data[645] = 6'b000110;
    assign data[646] = 6'b000110;
    assign data[647] = 6'b000111;
    assign data[648] = 6'b000111;
    assign data[649] = 6'b001000;
    assign data[650] = 6'b001000;
    assign data[651] = 6'b001001;
    assign data[652] = 6'b001001;
    assign data[653] = 6'b001010;
    assign data[654] = 6'b001011;
    assign data[655] = 6'b001011;
    assign data[656] = 6'b001100;
    assign data[657] = 6'b001101;
    assign data[658] = 6'b001101;
    assign data[659] = 6'b001110;
    assign data[660] = 6'b001111;
    assign data[661] = 6'b001111;
    assign data[662] = 6'b010000;
    assign data[663] = 6'b010001;
    assign data[664] = 6'b010010;
    assign data[665] = 6'b010011;
    assign data[666] = 6'b010100;
    assign data[667] = 6'b010100;
    assign data[668] = 6'b010101;
    assign data[669] = 6'b010110;
    assign data[670] = 6'b010111;
    assign data[671] = 6'b011000;
    assign data[672] = 6'b011001;
    assign data[673] = 6'b011010;
    assign data[674] = 6'b011011;
    assign data[675] = 6'b000011;
    assign data[676] = 6'b000011;
    assign data[677] = 6'b000011;
    assign data[678] = 6'b000011;
    assign data[679] = 6'b000011;
    assign data[680] = 6'b000011;
    assign data[681] = 6'b000100;
    assign data[682] = 6'b000100;
    assign data[683] = 6'b000100;
    assign data[684] = 6'b000100;
    assign data[685] = 6'b000101;
    assign data[686] = 6'b000101;
    assign data[687] = 6'b000101;
    assign data[688] = 6'b000110;
    assign data[689] = 6'b000110;
    assign data[690] = 6'b000110;
    assign data[691] = 6'b000111;
    assign data[692] = 6'b000111;
    assign data[693] = 6'b001000;
    assign data[694] = 6'b001000;
    assign data[695] = 6'b001001;
    assign data[696] = 6'b001001;
    assign data[697] = 6'b001010;
    assign data[698] = 6'b001010;
    assign data[699] = 6'b001011;
    assign data[700] = 6'b001100;
    assign data[701] = 6'b001100;
    assign data[702] = 6'b001101;
    assign data[703] = 6'b001110;
    assign data[704] = 6'b001110;
    assign data[705] = 6'b001111;
    assign data[706] = 6'b010000;
    assign data[707] = 6'b010001;
    assign data[708] = 6'b010001;
    assign data[709] = 6'b010010;
    assign data[710] = 6'b010011;
    assign data[711] = 6'b010100;
    assign data[712] = 6'b010101;
    assign data[713] = 6'b010110;
    assign data[714] = 6'b010110;
    assign data[715] = 6'b010111;
    assign data[716] = 6'b011000;
    assign data[717] = 6'b011001;
    assign data[718] = 6'b011010;
    assign data[719] = 6'b011011;
    assign data[720] = 6'b000011;
    assign data[721] = 6'b000011;
    assign data[722] = 6'b000100;
    assign data[723] = 6'b000100;
    assign data[724] = 6'b000100;
    assign data[725] = 6'b000100;
    assign data[726] = 6'b000100;
    assign data[727] = 6'b000100;
    assign data[728] = 6'b000100;
    assign data[729] = 6'b000101;
    assign data[730] = 6'b000101;
    assign data[731] = 6'b000101;
    assign data[732] = 6'b000110;
    assign data[733] = 6'b000110;
    assign data[734] = 6'b000110;
    assign data[735] = 6'b000111;
    assign data[736] = 6'b000111;
    assign data[737] = 6'b001000;
    assign data[738] = 6'b001000;
    assign data[739] = 6'b001001;
    assign data[740] = 6'b001001;
    assign data[741] = 6'b001010;
    assign data[742] = 6'b001010;
    assign data[743] = 6'b001011;
    assign data[744] = 6'b001011;
    assign data[745] = 6'b001100;
    assign data[746] = 6'b001101;
    assign data[747] = 6'b001101;
    assign data[748] = 6'b001110;
    assign data[749] = 6'b001111;
    assign data[750] = 6'b001111;
    assign data[751] = 6'b010000;
    assign data[752] = 6'b010001;
    assign data[753] = 6'b010010;
    assign data[754] = 6'b010011;
    assign data[755] = 6'b010011;
    assign data[756] = 6'b010100;
    assign data[757] = 6'b010101;
    assign data[758] = 6'b010110;
    assign data[759] = 6'b010111;
    assign data[760] = 6'b011000;
    assign data[761] = 6'b011001;
    assign data[762] = 6'b011010;
    assign data[763] = 6'b011010;
    assign data[764] = 6'b011011;
    assign data[765] = 6'b000100;
    assign data[766] = 6'b000100;
    assign data[767] = 6'b000100;
    assign data[768] = 6'b000100;
    assign data[769] = 6'b000100;
    assign data[770] = 6'b000100;
    assign data[771] = 6'b000100;
    assign data[772] = 6'b000101;
    assign data[773] = 6'b000101;
    assign data[774] = 6'b000101;
    assign data[775] = 6'b000101;
    assign data[776] = 6'b000110;
    assign data[777] = 6'b000110;
    assign data[778] = 6'b000110;
    assign data[779] = 6'b000111;
    assign data[780] = 6'b000111;
    assign data[781] = 6'b001000;
    assign data[782] = 6'b001000;
    assign data[783] = 6'b001001;
    assign data[784] = 6'b001001;
    assign data[785] = 6'b001010;
    assign data[786] = 6'b001010;
    assign data[787] = 6'b001011;
    assign data[788] = 6'b001011;
    assign data[789] = 6'b001100;
    assign data[790] = 6'b001100;
    assign data[791] = 6'b001101;
    assign data[792] = 6'b001110;
    assign data[793] = 6'b001110;
    assign data[794] = 6'b001111;
    assign data[795] = 6'b010000;
    assign data[796] = 6'b010001;
    assign data[797] = 6'b010001;
    assign data[798] = 6'b010010;
    assign data[799] = 6'b010011;
    assign data[800] = 6'b010100;
    assign data[801] = 6'b010101;
    assign data[802] = 6'b010101;
    assign data[803] = 6'b010110;
    assign data[804] = 6'b010111;
    assign data[805] = 6'b011000;
    assign data[806] = 6'b011001;
    assign data[807] = 6'b011010;
    assign data[808] = 6'b011011;
    assign data[809] = 6'b011100;
    assign data[810] = 6'b000100;
    assign data[811] = 6'b000100;
    assign data[812] = 6'b000100;
    assign data[813] = 6'b000101;
    assign data[814] = 6'b000101;
    assign data[815] = 6'b000101;
    assign data[816] = 6'b000101;
    assign data[817] = 6'b000101;
    assign data[818] = 6'b000101;
    assign data[819] = 6'b000110;
    assign data[820] = 6'b000110;
    assign data[821] = 6'b000110;
    assign data[822] = 6'b000111;
    assign data[823] = 6'b000111;
    assign data[824] = 6'b000111;
    assign data[825] = 6'b001000;
    assign data[826] = 6'b001000;
    assign data[827] = 6'b001001;
    assign data[828] = 6'b001001;
    assign data[829] = 6'b001001;
    assign data[830] = 6'b001010;
    assign data[831] = 6'b001011;
    assign data[832] = 6'b001011;
    assign data[833] = 6'b001100;
    assign data[834] = 6'b001100;
    assign data[835] = 6'b001101;
    assign data[836] = 6'b001110;
    assign data[837] = 6'b001110;
    assign data[838] = 6'b001111;
    assign data[839] = 6'b010000;
    assign data[840] = 6'b010000;
    assign data[841] = 6'b010001;
    assign data[842] = 6'b010010;
    assign data[843] = 6'b010011;
    assign data[844] = 6'b010011;
    assign data[845] = 6'b010100;
    assign data[846] = 6'b010101;
    assign data[847] = 6'b010110;
    assign data[848] = 6'b010111;
    assign data[849] = 6'b011000;
    assign data[850] = 6'b011000;
    assign data[851] = 6'b011001;
    assign data[852] = 6'b011010;
    assign data[853] = 6'b011011;
    assign data[854] = 6'b011100;
    assign data[855] = 6'b000101;
    assign data[856] = 6'b000101;
    assign data[857] = 6'b000101;
    assign data[858] = 6'b000101;
    assign data[859] = 6'b000101;
    assign data[860] = 6'b000101;
    assign data[861] = 6'b000110;
    assign data[862] = 6'b000110;
    assign data[863] = 6'b000110;
    assign data[864] = 6'b000110;
    assign data[865] = 6'b000110;
    assign data[866] = 6'b000111;
    assign data[867] = 6'b000111;
    assign data[868] = 6'b000111;
    assign data[869] = 6'b001000;
    assign data[870] = 6'b001000;
    assign data[871] = 6'b001001;
    assign data[872] = 6'b001001;
    assign data[873] = 6'b001001;
    assign data[874] = 6'b001010;
    assign data[875] = 6'b001010;
    assign data[876] = 6'b001011;
    assign data[877] = 6'b001100;
    assign data[878] = 6'b001100;
    assign data[879] = 6'b001101;
    assign data[880] = 6'b001101;
    assign data[881] = 6'b001110;
    assign data[882] = 6'b001111;
    assign data[883] = 6'b001111;
    assign data[884] = 6'b010000;
    assign data[885] = 6'b010001;
    assign data[886] = 6'b010010;
    assign data[887] = 6'b010010;
    assign data[888] = 6'b010011;
    assign data[889] = 6'b010100;
    assign data[890] = 6'b010101;
    assign data[891] = 6'b010101;
    assign data[892] = 6'b010110;
    assign data[893] = 6'b010111;
    assign data[894] = 6'b011000;
    assign data[895] = 6'b011001;
    assign data[896] = 6'b011010;
    assign data[897] = 6'b011011;
    assign data[898] = 6'b011100;
    assign data[899] = 6'b011101;
    assign data[900] = 6'b000101;
    assign data[901] = 6'b000110;
    assign data[902] = 6'b000110;
    assign data[903] = 6'b000110;
    assign data[904] = 6'b000110;
    assign data[905] = 6'b000110;
    assign data[906] = 6'b000110;
    assign data[907] = 6'b000110;
    assign data[908] = 6'b000110;
    assign data[909] = 6'b000111;
    assign data[910] = 6'b000111;
    assign data[911] = 6'b000111;
    assign data[912] = 6'b001000;
    assign data[913] = 6'b001000;
    assign data[914] = 6'b001000;
    assign data[915] = 6'b001001;
    assign data[916] = 6'b001001;
    assign data[917] = 6'b001010;
    assign data[918] = 6'b001010;
    assign data[919] = 6'b001010;
    assign data[920] = 6'b001011;
    assign data[921] = 6'b001100;
    assign data[922] = 6'b001100;
    assign data[923] = 6'b001101;
    assign data[924] = 6'b001101;
    assign data[925] = 6'b001110;
    assign data[926] = 6'b001111;
    assign data[927] = 6'b001111;
    assign data[928] = 6'b010000;
    assign data[929] = 6'b010001;
    assign data[930] = 6'b010001;
    assign data[931] = 6'b010010;
    assign data[932] = 6'b010011;
    assign data[933] = 6'b010100;
    assign data[934] = 6'b010100;
    assign data[935] = 6'b010101;
    assign data[936] = 6'b010110;
    assign data[937] = 6'b010111;
    assign data[938] = 6'b011000;
    assign data[939] = 6'b011000;
    assign data[940] = 6'b011001;
    assign data[941] = 6'b011010;
    assign data[942] = 6'b011011;
    assign data[943] = 6'b011100;
    assign data[944] = 6'b011101;
    assign data[945] = 6'b000110;
    assign data[946] = 6'b000110;
    assign data[947] = 6'b000110;
    assign data[948] = 6'b000110;
    assign data[949] = 6'b000110;
    assign data[950] = 6'b000110;
    assign data[951] = 6'b000111;
    assign data[952] = 6'b000111;
    assign data[953] = 6'b000111;
    assign data[954] = 6'b000111;
    assign data[955] = 6'b001000;
    assign data[956] = 6'b001000;
    assign data[957] = 6'b001000;
    assign data[958] = 6'b001000;
    assign data[959] = 6'b001001;
    assign data[960] = 6'b001001;
    assign data[961] = 6'b001010;
    assign data[962] = 6'b001010;
    assign data[963] = 6'b001011;
    assign data[964] = 6'b001011;
    assign data[965] = 6'b001100;
    assign data[966] = 6'b001100;
    assign data[967] = 6'b001101;
    assign data[968] = 6'b001101;
    assign data[969] = 6'b001110;
    assign data[970] = 6'b001110;
    assign data[971] = 6'b001111;
    assign data[972] = 6'b010000;
    assign data[973] = 6'b010000;
    assign data[974] = 6'b010001;
    assign data[975] = 6'b010010;
    assign data[976] = 6'b010010;
    assign data[977] = 6'b010011;
    assign data[978] = 6'b010100;
    assign data[979] = 6'b010101;
    assign data[980] = 6'b010110;
    assign data[981] = 6'b010110;
    assign data[982] = 6'b010111;
    assign data[983] = 6'b011000;
    assign data[984] = 6'b011001;
    assign data[985] = 6'b011010;
    assign data[986] = 6'b011011;
    assign data[987] = 6'b011100;
    assign data[988] = 6'b011100;
    assign data[989] = 6'b011101;
    assign data[990] = 6'b000111;
    assign data[991] = 6'b000111;
    assign data[992] = 6'b000111;
    assign data[993] = 6'b000111;
    assign data[994] = 6'b000111;
    assign data[995] = 6'b000111;
    assign data[996] = 6'b000111;
    assign data[997] = 6'b000111;
    assign data[998] = 6'b001000;
    assign data[999] = 6'b001000;
    assign data[1000] = 6'b001000;
    assign data[1001] = 6'b001000;
    assign data[1002] = 6'b001001;
    assign data[1003] = 6'b001001;
    assign data[1004] = 6'b001001;
    assign data[1005] = 6'b001010;
    assign data[1006] = 6'b001010;
    assign data[1007] = 6'b001011;
    assign data[1008] = 6'b001011;
    assign data[1009] = 6'b001100;
    assign data[1010] = 6'b001100;
    assign data[1011] = 6'b001101;
    assign data[1012] = 6'b001101;
    assign data[1013] = 6'b001110;
    assign data[1014] = 6'b001110;
    assign data[1015] = 6'b001111;
    assign data[1016] = 6'b010000;
    assign data[1017] = 6'b010000;
    assign data[1018] = 6'b010001;
    assign data[1019] = 6'b010010;
    assign data[1020] = 6'b010010;
    assign data[1021] = 6'b010011;
    assign data[1022] = 6'b010100;
    assign data[1023] = 6'b010100;
    assign data[1024] = 6'b010101;
    assign data[1025] = 6'b010110;
    assign data[1026] = 6'b010111;
    assign data[1027] = 6'b011000;
    assign data[1028] = 6'b011001;
    assign data[1029] = 6'b011001;
    assign data[1030] = 6'b011010;
    assign data[1031] = 6'b011011;
    assign data[1032] = 6'b011100;
    assign data[1033] = 6'b011101;
    assign data[1034] = 6'b011110;
    assign data[1035] = 6'b000111;
    assign data[1036] = 6'b000111;
    assign data[1037] = 6'b000111;
    assign data[1038] = 6'b000111;
    assign data[1039] = 6'b001000;
    assign data[1040] = 6'b001000;
    assign data[1041] = 6'b001000;
    assign data[1042] = 6'b001000;
    assign data[1043] = 6'b001000;
    assign data[1044] = 6'b001000;
    assign data[1045] = 6'b001001;
    assign data[1046] = 6'b001001;
    assign data[1047] = 6'b001001;
    assign data[1048] = 6'b001010;
    assign data[1049] = 6'b001010;
    assign data[1050] = 6'b001010;
    assign data[1051] = 6'b001011;
    assign data[1052] = 6'b001011;
    assign data[1053] = 6'b001100;
    assign data[1054] = 6'b001100;
    assign data[1055] = 6'b001101;
    assign data[1056] = 6'b001101;
    assign data[1057] = 6'b001110;
    assign data[1058] = 6'b001110;
    assign data[1059] = 6'b001111;
    assign data[1060] = 6'b001111;
    assign data[1061] = 6'b010000;
    assign data[1062] = 6'b010001;
    assign data[1063] = 6'b010001;
    assign data[1064] = 6'b010010;
    assign data[1065] = 6'b010011;
    assign data[1066] = 6'b010100;
    assign data[1067] = 6'b010100;
    assign data[1068] = 6'b010101;
    assign data[1069] = 6'b010110;
    assign data[1070] = 6'b010111;
    assign data[1071] = 6'b010111;
    assign data[1072] = 6'b011000;
    assign data[1073] = 6'b011001;
    assign data[1074] = 6'b011010;
    assign data[1075] = 6'b011011;
    assign data[1076] = 6'b011100;
    assign data[1077] = 6'b011101;
    assign data[1078] = 6'b011101;
    assign data[1079] = 6'b011110;
    assign data[1080] = 6'b001000;
    assign data[1081] = 6'b001000;
    assign data[1082] = 6'b001000;
    assign data[1083] = 6'b001000;
    assign data[1084] = 6'b001000;
    assign data[1085] = 6'b001000;
    assign data[1086] = 6'b001000;
    assign data[1087] = 6'b001001;
    assign data[1088] = 6'b001001;
    assign data[1089] = 6'b001001;
    assign data[1090] = 6'b001001;
    assign data[1091] = 6'b001010;
    assign data[1092] = 6'b001010;
    assign data[1093] = 6'b001010;
    assign data[1094] = 6'b001011;
    assign data[1095] = 6'b001011;
    assign data[1096] = 6'b001011;
    assign data[1097] = 6'b001100;
    assign data[1098] = 6'b001100;
    assign data[1099] = 6'b001101;
    assign data[1100] = 6'b001101;
    assign data[1101] = 6'b001110;
    assign data[1102] = 6'b001110;
    assign data[1103] = 6'b001111;
    assign data[1104] = 6'b001111;
    assign data[1105] = 6'b010000;
    assign data[1106] = 6'b010001;
    assign data[1107] = 6'b010001;
    assign data[1108] = 6'b010010;
    assign data[1109] = 6'b010011;
    assign data[1110] = 6'b010011;
    assign data[1111] = 6'b010100;
    assign data[1112] = 6'b010101;
    assign data[1113] = 6'b010110;
    assign data[1114] = 6'b010110;
    assign data[1115] = 6'b010111;
    assign data[1116] = 6'b011000;
    assign data[1117] = 6'b011001;
    assign data[1118] = 6'b011010;
    assign data[1119] = 6'b011010;
    assign data[1120] = 6'b011011;
    assign data[1121] = 6'b011100;
    assign data[1122] = 6'b011101;
    assign data[1123] = 6'b011110;
    assign data[1124] = 6'b011111;
    assign data[1125] = 6'b001001;
    assign data[1126] = 6'b001001;
    assign data[1127] = 6'b001001;
    assign data[1128] = 6'b001001;
    assign data[1129] = 6'b001001;
    assign data[1130] = 6'b001001;
    assign data[1131] = 6'b001001;
    assign data[1132] = 6'b001001;
    assign data[1133] = 6'b001001;
    assign data[1134] = 6'b001010;
    assign data[1135] = 6'b001010;
    assign data[1136] = 6'b001010;
    assign data[1137] = 6'b001011;
    assign data[1138] = 6'b001011;
    assign data[1139] = 6'b001011;
    assign data[1140] = 6'b001100;
    assign data[1141] = 6'b001100;
    assign data[1142] = 6'b001100;
    assign data[1143] = 6'b001101;
    assign data[1144] = 6'b001101;
    assign data[1145] = 6'b001110;
    assign data[1146] = 6'b001110;
    assign data[1147] = 6'b001111;
    assign data[1148] = 6'b001111;
    assign data[1149] = 6'b010000;
    assign data[1150] = 6'b010001;
    assign data[1151] = 6'b010001;
    assign data[1152] = 6'b010010;
    assign data[1153] = 6'b010011;
    assign data[1154] = 6'b010011;
    assign data[1155] = 6'b010100;
    assign data[1156] = 6'b010101;
    assign data[1157] = 6'b010101;
    assign data[1158] = 6'b010110;
    assign data[1159] = 6'b010111;
    assign data[1160] = 6'b011000;
    assign data[1161] = 6'b011000;
    assign data[1162] = 6'b011001;
    assign data[1163] = 6'b011010;
    assign data[1164] = 6'b011011;
    assign data[1165] = 6'b011100;
    assign data[1166] = 6'b011101;
    assign data[1167] = 6'b011110;
    assign data[1168] = 6'b011110;
    assign data[1169] = 6'b011111;
    assign data[1170] = 6'b001001;
    assign data[1171] = 6'b001001;
    assign data[1172] = 6'b001001;
    assign data[1173] = 6'b001001;
    assign data[1174] = 6'b001001;
    assign data[1175] = 6'b001010;
    assign data[1176] = 6'b001010;
    assign data[1177] = 6'b001010;
    assign data[1178] = 6'b001010;
    assign data[1179] = 6'b001010;
    assign data[1180] = 6'b001011;
    assign data[1181] = 6'b001011;
    assign data[1182] = 6'b001011;
    assign data[1183] = 6'b001100;
    assign data[1184] = 6'b001100;
    assign data[1185] = 6'b001100;
    assign data[1186] = 6'b001101;
    assign data[1187] = 6'b001101;
    assign data[1188] = 6'b001110;
    assign data[1189] = 6'b001110;
    assign data[1190] = 6'b001111;
    assign data[1191] = 6'b001111;
    assign data[1192] = 6'b010000;
    assign data[1193] = 6'b010000;
    assign data[1194] = 6'b010001;
    assign data[1195] = 6'b010001;
    assign data[1196] = 6'b010010;
    assign data[1197] = 6'b010011;
    assign data[1198] = 6'b010011;
    assign data[1199] = 6'b010100;
    assign data[1200] = 6'b010101;
    assign data[1201] = 6'b010101;
    assign data[1202] = 6'b010110;
    assign data[1203] = 6'b010111;
    assign data[1204] = 6'b010111;
    assign data[1205] = 6'b011000;
    assign data[1206] = 6'b011001;
    assign data[1207] = 6'b011010;
    assign data[1208] = 6'b011011;
    assign data[1209] = 6'b011011;
    assign data[1210] = 6'b011100;
    assign data[1211] = 6'b011101;
    assign data[1212] = 6'b011110;
    assign data[1213] = 6'b011111;
    assign data[1214] = 6'b100000;
    assign data[1215] = 6'b001010;
    assign data[1216] = 6'b001010;
    assign data[1217] = 6'b001010;
    assign data[1218] = 6'b001010;
    assign data[1219] = 6'b001010;
    assign data[1220] = 6'b001010;
    assign data[1221] = 6'b001010;
    assign data[1222] = 6'b001011;
    assign data[1223] = 6'b001011;
    assign data[1224] = 6'b001011;
    assign data[1225] = 6'b001011;
    assign data[1226] = 6'b001100;
    assign data[1227] = 6'b001100;
    assign data[1228] = 6'b001100;
    assign data[1229] = 6'b001101;
    assign data[1230] = 6'b001101;
    assign data[1231] = 6'b001101;
    assign data[1232] = 6'b001110;
    assign data[1233] = 6'b001110;
    assign data[1234] = 6'b001111;
    assign data[1235] = 6'b001111;
    assign data[1236] = 6'b010000;
    assign data[1237] = 6'b010000;
    assign data[1238] = 6'b010001;
    assign data[1239] = 6'b010001;
    assign data[1240] = 6'b010010;
    assign data[1241] = 6'b010011;
    assign data[1242] = 6'b010011;
    assign data[1243] = 6'b010100;
    assign data[1244] = 6'b010100;
    assign data[1245] = 6'b010101;
    assign data[1246] = 6'b010110;
    assign data[1247] = 6'b010111;
    assign data[1248] = 6'b010111;
    assign data[1249] = 6'b011000;
    assign data[1250] = 6'b011001;
    assign data[1251] = 6'b011010;
    assign data[1252] = 6'b011010;
    assign data[1253] = 6'b011011;
    assign data[1254] = 6'b011100;
    assign data[1255] = 6'b011101;
    assign data[1256] = 6'b011110;
    assign data[1257] = 6'b011111;
    assign data[1258] = 6'b100000;
    assign data[1259] = 6'b100000;
    assign data[1260] = 6'b001011;
    assign data[1261] = 6'b001011;
    assign data[1262] = 6'b001011;
    assign data[1263] = 6'b001011;
    assign data[1264] = 6'b001011;
    assign data[1265] = 6'b001011;
    assign data[1266] = 6'b001011;
    assign data[1267] = 6'b001011;
    assign data[1268] = 6'b001100;
    assign data[1269] = 6'b001100;
    assign data[1270] = 6'b001100;
    assign data[1271] = 6'b001100;
    assign data[1272] = 6'b001101;
    assign data[1273] = 6'b001101;
    assign data[1274] = 6'b001101;
    assign data[1275] = 6'b001110;
    assign data[1276] = 6'b001110;
    assign data[1277] = 6'b001110;
    assign data[1278] = 6'b001111;
    assign data[1279] = 6'b001111;
    assign data[1280] = 6'b010000;
    assign data[1281] = 6'b010000;
    assign data[1282] = 6'b010001;
    assign data[1283] = 6'b010001;
    assign data[1284] = 6'b010010;
    assign data[1285] = 6'b010011;
    assign data[1286] = 6'b010011;
    assign data[1287] = 6'b010100;
    assign data[1288] = 6'b010100;
    assign data[1289] = 6'b010101;
    assign data[1290] = 6'b010110;
    assign data[1291] = 6'b010110;
    assign data[1292] = 6'b010111;
    assign data[1293] = 6'b011000;
    assign data[1294] = 6'b011001;
    assign data[1295] = 6'b011001;
    assign data[1296] = 6'b011010;
    assign data[1297] = 6'b011011;
    assign data[1298] = 6'b011100;
    assign data[1299] = 6'b011101;
    assign data[1300] = 6'b011101;
    assign data[1301] = 6'b011110;
    assign data[1302] = 6'b011111;
    assign data[1303] = 6'b100000;
    assign data[1304] = 6'b100001;
    assign data[1305] = 6'b001011;
    assign data[1306] = 6'b001011;
    assign data[1307] = 6'b001011;
    assign data[1308] = 6'b001100;
    assign data[1309] = 6'b001100;
    assign data[1310] = 6'b001100;
    assign data[1311] = 6'b001100;
    assign data[1312] = 6'b001100;
    assign data[1313] = 6'b001100;
    assign data[1314] = 6'b001101;
    assign data[1315] = 6'b001101;
    assign data[1316] = 6'b001101;
    assign data[1317] = 6'b001101;
    assign data[1318] = 6'b001110;
    assign data[1319] = 6'b001110;
    assign data[1320] = 6'b001110;
    assign data[1321] = 6'b001111;
    assign data[1322] = 6'b001111;
    assign data[1323] = 6'b010000;
    assign data[1324] = 6'b010000;
    assign data[1325] = 6'b010001;
    assign data[1326] = 6'b010001;
    assign data[1327] = 6'b010010;
    assign data[1328] = 6'b010010;
    assign data[1329] = 6'b010011;
    assign data[1330] = 6'b010011;
    assign data[1331] = 6'b010100;
    assign data[1332] = 6'b010100;
    assign data[1333] = 6'b010101;
    assign data[1334] = 6'b010110;
    assign data[1335] = 6'b010110;
    assign data[1336] = 6'b010111;
    assign data[1337] = 6'b011000;
    assign data[1338] = 6'b011001;
    assign data[1339] = 6'b011001;
    assign data[1340] = 6'b011010;
    assign data[1341] = 6'b011011;
    assign data[1342] = 6'b011100;
    assign data[1343] = 6'b011100;
    assign data[1344] = 6'b011101;
    assign data[1345] = 6'b011110;
    assign data[1346] = 6'b011111;
    assign data[1347] = 6'b100000;
    assign data[1348] = 6'b100001;
    assign data[1349] = 6'b100010;
    assign data[1350] = 6'b001100;
    assign data[1351] = 6'b001100;
    assign data[1352] = 6'b001100;
    assign data[1353] = 6'b001100;
    assign data[1354] = 6'b001100;
    assign data[1355] = 6'b001101;
    assign data[1356] = 6'b001101;
    assign data[1357] = 6'b001101;
    assign data[1358] = 6'b001101;
    assign data[1359] = 6'b001101;
    assign data[1360] = 6'b001110;
    assign data[1361] = 6'b001110;
    assign data[1362] = 6'b001110;
    assign data[1363] = 6'b001110;
    assign data[1364] = 6'b001111;
    assign data[1365] = 6'b001111;
    assign data[1366] = 6'b001111;
    assign data[1367] = 6'b010000;
    assign data[1368] = 6'b010000;
    assign data[1369] = 6'b010001;
    assign data[1370] = 6'b010001;
    assign data[1371] = 6'b010010;
    assign data[1372] = 6'b010010;
    assign data[1373] = 6'b010011;
    assign data[1374] = 6'b010011;
    assign data[1375] = 6'b010100;
    assign data[1376] = 6'b010101;
    assign data[1377] = 6'b010101;
    assign data[1378] = 6'b010110;
    assign data[1379] = 6'b010110;
    assign data[1380] = 6'b010111;
    assign data[1381] = 6'b011000;
    assign data[1382] = 6'b011001;
    assign data[1383] = 6'b011001;
    assign data[1384] = 6'b011010;
    assign data[1385] = 6'b011011;
    assign data[1386] = 6'b011011;
    assign data[1387] = 6'b011100;
    assign data[1388] = 6'b011101;
    assign data[1389] = 6'b011110;
    assign data[1390] = 6'b011111;
    assign data[1391] = 6'b100000;
    assign data[1392] = 6'b100000;
    assign data[1393] = 6'b100001;
    assign data[1394] = 6'b100010;
    assign data[1395] = 6'b001101;
    assign data[1396] = 6'b001101;
    assign data[1397] = 6'b001101;
    assign data[1398] = 6'b001101;
    assign data[1399] = 6'b001101;
    assign data[1400] = 6'b001101;
    assign data[1401] = 6'b001101;
    assign data[1402] = 6'b001110;
    assign data[1403] = 6'b001110;
    assign data[1404] = 6'b001110;
    assign data[1405] = 6'b001110;
    assign data[1406] = 6'b001111;
    assign data[1407] = 6'b001111;
    assign data[1408] = 6'b001111;
    assign data[1409] = 6'b001111;
    assign data[1410] = 6'b010000;
    assign data[1411] = 6'b010000;
    assign data[1412] = 6'b010001;
    assign data[1413] = 6'b010001;
    assign data[1414] = 6'b010010;
    assign data[1415] = 6'b010010;
    assign data[1416] = 6'b010010;
    assign data[1417] = 6'b010011;
    assign data[1418] = 6'b010100;
    assign data[1419] = 6'b010100;
    assign data[1420] = 6'b010101;
    assign data[1421] = 6'b010101;
    assign data[1422] = 6'b010110;
    assign data[1423] = 6'b010110;
    assign data[1424] = 6'b010111;
    assign data[1425] = 6'b011000;
    assign data[1426] = 6'b011000;
    assign data[1427] = 6'b011001;
    assign data[1428] = 6'b011010;
    assign data[1429] = 6'b011011;
    assign data[1430] = 6'b011011;
    assign data[1431] = 6'b011100;
    assign data[1432] = 6'b011101;
    assign data[1433] = 6'b011110;
    assign data[1434] = 6'b011111;
    assign data[1435] = 6'b011111;
    assign data[1436] = 6'b100000;
    assign data[1437] = 6'b100001;
    assign data[1438] = 6'b100010;
    assign data[1439] = 6'b100011;
    assign data[1440] = 6'b001110;
    assign data[1441] = 6'b001110;
    assign data[1442] = 6'b001110;
    assign data[1443] = 6'b001110;
    assign data[1444] = 6'b001110;
    assign data[1445] = 6'b001110;
    assign data[1446] = 6'b001110;
    assign data[1447] = 6'b001110;
    assign data[1448] = 6'b001111;
    assign data[1449] = 6'b001111;
    assign data[1450] = 6'b001111;
    assign data[1451] = 6'b001111;
    assign data[1452] = 6'b010000;
    assign data[1453] = 6'b010000;
    assign data[1454] = 6'b010000;
    assign data[1455] = 6'b010001;
    assign data[1456] = 6'b010001;
    assign data[1457] = 6'b010001;
    assign data[1458] = 6'b010010;
    assign data[1459] = 6'b010010;
    assign data[1460] = 6'b010011;
    assign data[1461] = 6'b010011;
    assign data[1462] = 6'b010100;
    assign data[1463] = 6'b010100;
    assign data[1464] = 6'b010101;
    assign data[1465] = 6'b010101;
    assign data[1466] = 6'b010110;
    assign data[1467] = 6'b010111;
    assign data[1468] = 6'b010111;
    assign data[1469] = 6'b011000;
    assign data[1470] = 6'b011001;
    assign data[1471] = 6'b011001;
    assign data[1472] = 6'b011010;
    assign data[1473] = 6'b011011;
    assign data[1474] = 6'b011011;
    assign data[1475] = 6'b011100;
    assign data[1476] = 6'b011101;
    assign data[1477] = 6'b011110;
    assign data[1478] = 6'b011110;
    assign data[1479] = 6'b011111;
    assign data[1480] = 6'b100000;
    assign data[1481] = 6'b100001;
    assign data[1482] = 6'b100010;
    assign data[1483] = 6'b100011;
    assign data[1484] = 6'b100011;
    assign data[1485] = 6'b001111;
    assign data[1486] = 6'b001111;
    assign data[1487] = 6'b001111;
    assign data[1488] = 6'b001111;
    assign data[1489] = 6'b001111;
    assign data[1490] = 6'b001111;
    assign data[1491] = 6'b001111;
    assign data[1492] = 6'b001111;
    assign data[1493] = 6'b001111;
    assign data[1494] = 6'b010000;
    assign data[1495] = 6'b010000;
    assign data[1496] = 6'b010000;
    assign data[1497] = 6'b010000;
    assign data[1498] = 6'b010001;
    assign data[1499] = 6'b010001;
    assign data[1500] = 6'b010001;
    assign data[1501] = 6'b010010;
    assign data[1502] = 6'b010010;
    assign data[1503] = 6'b010011;
    assign data[1504] = 6'b010011;
    assign data[1505] = 6'b010100;
    assign data[1506] = 6'b010100;
    assign data[1507] = 6'b010100;
    assign data[1508] = 6'b010101;
    assign data[1509] = 6'b010110;
    assign data[1510] = 6'b010110;
    assign data[1511] = 6'b010111;
    assign data[1512] = 6'b010111;
    assign data[1513] = 6'b011000;
    assign data[1514] = 6'b011001;
    assign data[1515] = 6'b011001;
    assign data[1516] = 6'b011010;
    assign data[1517] = 6'b011011;
    assign data[1518] = 6'b011011;
    assign data[1519] = 6'b011100;
    assign data[1520] = 6'b011101;
    assign data[1521] = 6'b011110;
    assign data[1522] = 6'b011110;
    assign data[1523] = 6'b011111;
    assign data[1524] = 6'b100000;
    assign data[1525] = 6'b100001;
    assign data[1526] = 6'b100010;
    assign data[1527] = 6'b100010;
    assign data[1528] = 6'b100011;
    assign data[1529] = 6'b100100;
    assign data[1530] = 6'b001111;
    assign data[1531] = 6'b001111;
    assign data[1532] = 6'b001111;
    assign data[1533] = 6'b001111;
    assign data[1534] = 6'b010000;
    assign data[1535] = 6'b010000;
    assign data[1536] = 6'b010000;
    assign data[1537] = 6'b010000;
    assign data[1538] = 6'b010000;
    assign data[1539] = 6'b010000;
    assign data[1540] = 6'b010001;
    assign data[1541] = 6'b010001;
    assign data[1542] = 6'b010001;
    assign data[1543] = 6'b010010;
    assign data[1544] = 6'b010010;
    assign data[1545] = 6'b010010;
    assign data[1546] = 6'b010011;
    assign data[1547] = 6'b010011;
    assign data[1548] = 6'b010011;
    assign data[1549] = 6'b010100;
    assign data[1550] = 6'b010100;
    assign data[1551] = 6'b010101;
    assign data[1552] = 6'b010101;
    assign data[1553] = 6'b010110;
    assign data[1554] = 6'b010110;
    assign data[1555] = 6'b010111;
    assign data[1556] = 6'b010111;
    assign data[1557] = 6'b011000;
    assign data[1558] = 6'b011001;
    assign data[1559] = 6'b011001;
    assign data[1560] = 6'b011010;
    assign data[1561] = 6'b011011;
    assign data[1562] = 6'b011011;
    assign data[1563] = 6'b011100;
    assign data[1564] = 6'b011101;
    assign data[1565] = 6'b011101;
    assign data[1566] = 6'b011110;
    assign data[1567] = 6'b011111;
    assign data[1568] = 6'b100000;
    assign data[1569] = 6'b100001;
    assign data[1570] = 6'b100001;
    assign data[1571] = 6'b100010;
    assign data[1572] = 6'b100011;
    assign data[1573] = 6'b100100;
    assign data[1574] = 6'b100101;
    assign data[1575] = 6'b010000;
    assign data[1576] = 6'b010000;
    assign data[1577] = 6'b010000;
    assign data[1578] = 6'b010000;
    assign data[1579] = 6'b010000;
    assign data[1580] = 6'b010001;
    assign data[1581] = 6'b010001;
    assign data[1582] = 6'b010001;
    assign data[1583] = 6'b010001;
    assign data[1584] = 6'b010001;
    assign data[1585] = 6'b010001;
    assign data[1586] = 6'b010010;
    assign data[1587] = 6'b010010;
    assign data[1588] = 6'b010010;
    assign data[1589] = 6'b010011;
    assign data[1590] = 6'b010011;
    assign data[1591] = 6'b010011;
    assign data[1592] = 6'b010100;
    assign data[1593] = 6'b010100;
    assign data[1594] = 6'b010101;
    assign data[1595] = 6'b010101;
    assign data[1596] = 6'b010110;
    assign data[1597] = 6'b010110;
    assign data[1598] = 6'b010111;
    assign data[1599] = 6'b010111;
    assign data[1600] = 6'b011000;
    assign data[1601] = 6'b011000;
    assign data[1602] = 6'b011001;
    assign data[1603] = 6'b011001;
    assign data[1604] = 6'b011010;
    assign data[1605] = 6'b011011;
    assign data[1606] = 6'b011011;
    assign data[1607] = 6'b011100;
    assign data[1608] = 6'b011101;
    assign data[1609] = 6'b011101;
    assign data[1610] = 6'b011110;
    assign data[1611] = 6'b011111;
    assign data[1612] = 6'b100000;
    assign data[1613] = 6'b100000;
    assign data[1614] = 6'b100001;
    assign data[1615] = 6'b100010;
    assign data[1616] = 6'b100011;
    assign data[1617] = 6'b100100;
    assign data[1618] = 6'b100101;
    assign data[1619] = 6'b100101;
    assign data[1620] = 6'b010001;
    assign data[1621] = 6'b010001;
    assign data[1622] = 6'b010001;
    assign data[1623] = 6'b010001;
    assign data[1624] = 6'b010001;
    assign data[1625] = 6'b010001;
    assign data[1626] = 6'b010010;
    assign data[1627] = 6'b010010;
    assign data[1628] = 6'b010010;
    assign data[1629] = 6'b010010;
    assign data[1630] = 6'b010010;
    assign data[1631] = 6'b010011;
    assign data[1632] = 6'b010011;
    assign data[1633] = 6'b010011;
    assign data[1634] = 6'b010100;
    assign data[1635] = 6'b010100;
    assign data[1636] = 6'b010100;
    assign data[1637] = 6'b010101;
    assign data[1638] = 6'b010101;
    assign data[1639] = 6'b010101;
    assign data[1640] = 6'b010110;
    assign data[1641] = 6'b010110;
    assign data[1642] = 6'b010111;
    assign data[1643] = 6'b010111;
    assign data[1644] = 6'b011000;
    assign data[1645] = 6'b011000;
    assign data[1646] = 6'b011001;
    assign data[1647] = 6'b011010;
    assign data[1648] = 6'b011010;
    assign data[1649] = 6'b011011;
    assign data[1650] = 6'b011011;
    assign data[1651] = 6'b011100;
    assign data[1652] = 6'b011101;
    assign data[1653] = 6'b011110;
    assign data[1654] = 6'b011110;
    assign data[1655] = 6'b011111;
    assign data[1656] = 6'b100000;
    assign data[1657] = 6'b100000;
    assign data[1658] = 6'b100001;
    assign data[1659] = 6'b100010;
    assign data[1660] = 6'b100011;
    assign data[1661] = 6'b100100;
    assign data[1662] = 6'b100100;
    assign data[1663] = 6'b100101;
    assign data[1664] = 6'b100110;
    assign data[1665] = 6'b010010;
    assign data[1666] = 6'b010010;
    assign data[1667] = 6'b010010;
    assign data[1668] = 6'b010010;
    assign data[1669] = 6'b010010;
    assign data[1670] = 6'b010010;
    assign data[1671] = 6'b010010;
    assign data[1672] = 6'b010011;
    assign data[1673] = 6'b010011;
    assign data[1674] = 6'b010011;
    assign data[1675] = 6'b010011;
    assign data[1676] = 6'b010011;
    assign data[1677] = 6'b010100;
    assign data[1678] = 6'b010100;
    assign data[1679] = 6'b010100;
    assign data[1680] = 6'b010101;
    assign data[1681] = 6'b010101;
    assign data[1682] = 6'b010101;
    assign data[1683] = 6'b010110;
    assign data[1684] = 6'b010110;
    assign data[1685] = 6'b010111;
    assign data[1686] = 6'b010111;
    assign data[1687] = 6'b011000;
    assign data[1688] = 6'b011000;
    assign data[1689] = 6'b011001;
    assign data[1690] = 6'b011001;
    assign data[1691] = 6'b011010;
    assign data[1692] = 6'b011010;
    assign data[1693] = 6'b011011;
    assign data[1694] = 6'b011100;
    assign data[1695] = 6'b011100;
    assign data[1696] = 6'b011101;
    assign data[1697] = 6'b011110;
    assign data[1698] = 6'b011110;
    assign data[1699] = 6'b011111;
    assign data[1700] = 6'b100000;
    assign data[1701] = 6'b100000;
    assign data[1702] = 6'b100001;
    assign data[1703] = 6'b100010;
    assign data[1704] = 6'b100011;
    assign data[1705] = 6'b100100;
    assign data[1706] = 6'b100100;
    assign data[1707] = 6'b100101;
    assign data[1708] = 6'b100110;
    assign data[1709] = 6'b100111;
    assign data[1710] = 6'b010011;
    assign data[1711] = 6'b010011;
    assign data[1712] = 6'b010011;
    assign data[1713] = 6'b010011;
    assign data[1714] = 6'b010011;
    assign data[1715] = 6'b010011;
    assign data[1716] = 6'b010011;
    assign data[1717] = 6'b010011;
    assign data[1718] = 6'b010100;
    assign data[1719] = 6'b010100;
    assign data[1720] = 6'b010100;
    assign data[1721] = 6'b010100;
    assign data[1722] = 6'b010101;
    assign data[1723] = 6'b010101;
    assign data[1724] = 6'b010101;
    assign data[1725] = 6'b010110;
    assign data[1726] = 6'b010110;
    assign data[1727] = 6'b010110;
    assign data[1728] = 6'b010111;
    assign data[1729] = 6'b010111;
    assign data[1730] = 6'b011000;
    assign data[1731] = 6'b011000;
    assign data[1732] = 6'b011001;
    assign data[1733] = 6'b011001;
    assign data[1734] = 6'b011010;
    assign data[1735] = 6'b011010;
    assign data[1736] = 6'b011011;
    assign data[1737] = 6'b011011;
    assign data[1738] = 6'b011100;
    assign data[1739] = 6'b011100;
    assign data[1740] = 6'b011101;
    assign data[1741] = 6'b011110;
    assign data[1742] = 6'b011110;
    assign data[1743] = 6'b011111;
    assign data[1744] = 6'b100000;
    assign data[1745] = 6'b100000;
    assign data[1746] = 6'b100001;
    assign data[1747] = 6'b100010;
    assign data[1748] = 6'b100011;
    assign data[1749] = 6'b100011;
    assign data[1750] = 6'b100100;
    assign data[1751] = 6'b100101;
    assign data[1752] = 6'b100110;
    assign data[1753] = 6'b100111;
    assign data[1754] = 6'b101000;
    assign data[1755] = 6'b010100;
    assign data[1756] = 6'b010100;
    assign data[1757] = 6'b010100;
    assign data[1758] = 6'b010100;
    assign data[1759] = 6'b010100;
    assign data[1760] = 6'b010100;
    assign data[1761] = 6'b010100;
    assign data[1762] = 6'b010100;
    assign data[1763] = 6'b010101;
    assign data[1764] = 6'b010101;
    assign data[1765] = 6'b010101;
    assign data[1766] = 6'b010101;
    assign data[1767] = 6'b010101;
    assign data[1768] = 6'b010110;
    assign data[1769] = 6'b010110;
    assign data[1770] = 6'b010110;
    assign data[1771] = 6'b010111;
    assign data[1772] = 6'b010111;
    assign data[1773] = 6'b011000;
    assign data[1774] = 6'b011000;
    assign data[1775] = 6'b011000;
    assign data[1776] = 6'b011001;
    assign data[1777] = 6'b011001;
    assign data[1778] = 6'b011010;
    assign data[1779] = 6'b011010;
    assign data[1780] = 6'b011011;
    assign data[1781] = 6'b011011;
    assign data[1782] = 6'b011100;
    assign data[1783] = 6'b011101;
    assign data[1784] = 6'b011101;
    assign data[1785] = 6'b011110;
    assign data[1786] = 6'b011111;
    assign data[1787] = 6'b011111;
    assign data[1788] = 6'b100000;
    assign data[1789] = 6'b100001;
    assign data[1790] = 6'b100001;
    assign data[1791] = 6'b100010;
    assign data[1792] = 6'b100011;
    assign data[1793] = 6'b100011;
    assign data[1794] = 6'b100100;
    assign data[1795] = 6'b100101;
    assign data[1796] = 6'b100110;
    assign data[1797] = 6'b100111;
    assign data[1798] = 6'b100111;
    assign data[1799] = 6'b101000;
    assign data[1800] = 6'b010101;
    assign data[1801] = 6'b010101;
    assign data[1802] = 6'b010101;
    assign data[1803] = 6'b010101;
    assign data[1804] = 6'b010101;
    assign data[1805] = 6'b010101;
    assign data[1806] = 6'b010101;
    assign data[1807] = 6'b010101;
    assign data[1808] = 6'b010101;
    assign data[1809] = 6'b010110;
    assign data[1810] = 6'b010110;
    assign data[1811] = 6'b010110;
    assign data[1812] = 6'b010110;
    assign data[1813] = 6'b010111;
    assign data[1814] = 6'b010111;
    assign data[1815] = 6'b010111;
    assign data[1816] = 6'b011000;
    assign data[1817] = 6'b011000;
    assign data[1818] = 6'b011000;
    assign data[1819] = 6'b011001;
    assign data[1820] = 6'b011001;
    assign data[1821] = 6'b011010;
    assign data[1822] = 6'b011010;
    assign data[1823] = 6'b011011;
    assign data[1824] = 6'b011011;
    assign data[1825] = 6'b011100;
    assign data[1826] = 6'b011100;
    assign data[1827] = 6'b011101;
    assign data[1828] = 6'b011101;
    assign data[1829] = 6'b011110;
    assign data[1830] = 6'b011111;
    assign data[1831] = 6'b011111;
    assign data[1832] = 6'b100000;
    assign data[1833] = 6'b100001;
    assign data[1834] = 6'b100001;
    assign data[1835] = 6'b100010;
    assign data[1836] = 6'b100011;
    assign data[1837] = 6'b100100;
    assign data[1838] = 6'b100100;
    assign data[1839] = 6'b100101;
    assign data[1840] = 6'b100110;
    assign data[1841] = 6'b100111;
    assign data[1842] = 6'b100111;
    assign data[1843] = 6'b101000;
    assign data[1844] = 6'b101001;
    assign data[1845] = 6'b010110;
    assign data[1846] = 6'b010110;
    assign data[1847] = 6'b010110;
    assign data[1848] = 6'b010110;
    assign data[1849] = 6'b010110;
    assign data[1850] = 6'b010110;
    assign data[1851] = 6'b010110;
    assign data[1852] = 6'b010110;
    assign data[1853] = 6'b010110;
    assign data[1854] = 6'b010111;
    assign data[1855] = 6'b010111;
    assign data[1856] = 6'b010111;
    assign data[1857] = 6'b010111;
    assign data[1858] = 6'b011000;
    assign data[1859] = 6'b011000;
    assign data[1860] = 6'b011000;
    assign data[1861] = 6'b011001;
    assign data[1862] = 6'b011001;
    assign data[1863] = 6'b011001;
    assign data[1864] = 6'b011010;
    assign data[1865] = 6'b011010;
    assign data[1866] = 6'b011011;
    assign data[1867] = 6'b011011;
    assign data[1868] = 6'b011100;
    assign data[1869] = 6'b011100;
    assign data[1870] = 6'b011101;
    assign data[1871] = 6'b011101;
    assign data[1872] = 6'b011110;
    assign data[1873] = 6'b011110;
    assign data[1874] = 6'b011111;
    assign data[1875] = 6'b100000;
    assign data[1876] = 6'b100000;
    assign data[1877] = 6'b100001;
    assign data[1878] = 6'b100010;
    assign data[1879] = 6'b100010;
    assign data[1880] = 6'b100011;
    assign data[1881] = 6'b100100;
    assign data[1882] = 6'b100100;
    assign data[1883] = 6'b100101;
    assign data[1884] = 6'b100110;
    assign data[1885] = 6'b100111;
    assign data[1886] = 6'b100111;
    assign data[1887] = 6'b101000;
    assign data[1888] = 6'b101001;
    assign data[1889] = 6'b101010;
    assign data[1890] = 6'b010111;
    assign data[1891] = 6'b010111;
    assign data[1892] = 6'b010111;
    assign data[1893] = 6'b010111;
    assign data[1894] = 6'b010111;
    assign data[1895] = 6'b010111;
    assign data[1896] = 6'b010111;
    assign data[1897] = 6'b010111;
    assign data[1898] = 6'b010111;
    assign data[1899] = 6'b011000;
    assign data[1900] = 6'b011000;
    assign data[1901] = 6'b011000;
    assign data[1902] = 6'b011000;
    assign data[1903] = 6'b011001;
    assign data[1904] = 6'b011001;
    assign data[1905] = 6'b011001;
    assign data[1906] = 6'b011010;
    assign data[1907] = 6'b011010;
    assign data[1908] = 6'b011010;
    assign data[1909] = 6'b011011;
    assign data[1910] = 6'b011011;
    assign data[1911] = 6'b011100;
    assign data[1912] = 6'b011100;
    assign data[1913] = 6'b011101;
    assign data[1914] = 6'b011101;
    assign data[1915] = 6'b011110;
    assign data[1916] = 6'b011110;
    assign data[1917] = 6'b011111;
    assign data[1918] = 6'b011111;
    assign data[1919] = 6'b100000;
    assign data[1920] = 6'b100000;
    assign data[1921] = 6'b100001;
    assign data[1922] = 6'b100010;
    assign data[1923] = 6'b100010;
    assign data[1924] = 6'b100011;
    assign data[1925] = 6'b100100;
    assign data[1926] = 6'b100100;
    assign data[1927] = 6'b100101;
    assign data[1928] = 6'b100110;
    assign data[1929] = 6'b100111;
    assign data[1930] = 6'b100111;
    assign data[1931] = 6'b101000;
    assign data[1932] = 6'b101001;
    assign data[1933] = 6'b101010;
    assign data[1934] = 6'b101011;
    assign data[1935] = 6'b010111;
    assign data[1936] = 6'b010111;
    assign data[1937] = 6'b011000;
    assign data[1938] = 6'b011000;
    assign data[1939] = 6'b011000;
    assign data[1940] = 6'b011000;
    assign data[1941] = 6'b011000;
    assign data[1942] = 6'b011000;
    assign data[1943] = 6'b011000;
    assign data[1944] = 6'b011000;
    assign data[1945] = 6'b011001;
    assign data[1946] = 6'b011001;
    assign data[1947] = 6'b011001;
    assign data[1948] = 6'b011001;
    assign data[1949] = 6'b011010;
    assign data[1950] = 6'b011010;
    assign data[1951] = 6'b011010;
    assign data[1952] = 6'b011011;
    assign data[1953] = 6'b011011;
    assign data[1954] = 6'b011100;
    assign data[1955] = 6'b011100;
    assign data[1956] = 6'b011100;
    assign data[1957] = 6'b011101;
    assign data[1958] = 6'b011101;
    assign data[1959] = 6'b011110;
    assign data[1960] = 6'b011110;
    assign data[1961] = 6'b011111;
    assign data[1962] = 6'b100000;
    assign data[1963] = 6'b100000;
    assign data[1964] = 6'b100001;
    assign data[1965] = 6'b100001;
    assign data[1966] = 6'b100010;
    assign data[1967] = 6'b100011;
    assign data[1968] = 6'b100011;
    assign data[1969] = 6'b100100;
    assign data[1970] = 6'b100101;
    assign data[1971] = 6'b100101;
    assign data[1972] = 6'b100110;
    assign data[1973] = 6'b100111;
    assign data[1974] = 6'b100111;
    assign data[1975] = 6'b101000;
    assign data[1976] = 6'b101001;
    assign data[1977] = 6'b101010;
    assign data[1978] = 6'b101011;
    assign data[1979] = 6'b101011;
    assign data[1980] = 6'b011000;
    assign data[1981] = 6'b011000;
    assign data[1982] = 6'b011001;
    assign data[1983] = 6'b011001;
    assign data[1984] = 6'b011001;
    assign data[1985] = 6'b011001;
    assign data[1986] = 6'b011001;
    assign data[1987] = 6'b011001;
    assign data[1988] = 6'b011001;
    assign data[1989] = 6'b011001;
    assign data[1990] = 6'b011010;
    assign data[1991] = 6'b011010;
    assign data[1992] = 6'b011010;
    assign data[1993] = 6'b011010;
    assign data[1994] = 6'b011011;
    assign data[1995] = 6'b011011;
    assign data[1996] = 6'b011011;
    assign data[1997] = 6'b011100;
    assign data[1998] = 6'b011100;
    assign data[1999] = 6'b011101;
    assign data[2000] = 6'b011101;
    assign data[2001] = 6'b011101;
    assign data[2002] = 6'b011110;
    assign data[2003] = 6'b011110;
    assign data[2004] = 6'b011111;
    assign data[2005] = 6'b011111;
    assign data[2006] = 6'b100000;
    assign data[2007] = 6'b100000;
    assign data[2008] = 6'b100001;
    assign data[2009] = 6'b100010;
    assign data[2010] = 6'b100010;
    assign data[2011] = 6'b100011;
    assign data[2012] = 6'b100011;
    assign data[2013] = 6'b100100;
    assign data[2014] = 6'b100101;
    assign data[2015] = 6'b100101;
    assign data[2016] = 6'b100110;
    assign data[2017] = 6'b100111;
    assign data[2018] = 6'b101000;
    assign data[2019] = 6'b101000;
    assign data[2020] = 6'b101001;
    assign data[2021] = 6'b101010;
    assign data[2022] = 6'b101011;
    assign data[2023] = 6'b101011;
    assign data[2024] = 6'b101100;
    assign data[2025] = 6'b011001;
    assign data[2026] = 6'b011001;
    assign data[2027] = 6'b011001;
    assign data[2028] = 6'b011010;
    assign data[2029] = 6'b011010;
    assign data[2030] = 6'b011010;
    assign data[2031] = 6'b011010;
    assign data[2032] = 6'b011010;
    assign data[2033] = 6'b011010;
    assign data[2034] = 6'b011010;
    assign data[2035] = 6'b011011;
    assign data[2036] = 6'b011011;
    assign data[2037] = 6'b011011;
    assign data[2038] = 6'b011011;
    assign data[2039] = 6'b011100;
    assign data[2040] = 6'b011100;
    assign data[2041] = 6'b011100;
    assign data[2042] = 6'b011101;
    assign data[2043] = 6'b011101;
    assign data[2044] = 6'b011101;
    assign data[2045] = 6'b011110;
    assign data[2046] = 6'b011110;
    assign data[2047] = 6'b011111;
    assign data[2048] = 6'b011111;
    assign data[2049] = 6'b100000;
    assign data[2050] = 6'b100000;
    assign data[2051] = 6'b100001;
    assign data[2052] = 6'b100001;
    assign data[2053] = 6'b100010;
    assign data[2054] = 6'b100010;
    assign data[2055] = 6'b100011;
    assign data[2056] = 6'b100100;
    assign data[2057] = 6'b100100;
    assign data[2058] = 6'b100101;
    assign data[2059] = 6'b100110;
    assign data[2060] = 6'b100110;
    assign data[2061] = 6'b100111;
    assign data[2062] = 6'b101000;
    assign data[2063] = 6'b101000;
    assign data[2064] = 6'b101001;
    assign data[2065] = 6'b101010;
    assign data[2066] = 6'b101011;
    assign data[2067] = 6'b101011;
    assign data[2068] = 6'b101100;
    assign data[2069] = 6'b101101;
    assign data[2070] = 6'b011010;
    assign data[2071] = 6'b011010;
    assign data[2072] = 6'b011010;
    assign data[2073] = 6'b011011;
    assign data[2074] = 6'b011011;
    assign data[2075] = 6'b011011;
    assign data[2076] = 6'b011011;
    assign data[2077] = 6'b011011;
    assign data[2078] = 6'b011011;
    assign data[2079] = 6'b011011;
    assign data[2080] = 6'b011100;
    assign data[2081] = 6'b011100;
    assign data[2082] = 6'b011100;
    assign data[2083] = 6'b011100;
    assign data[2084] = 6'b011101;
    assign data[2085] = 6'b011101;
    assign data[2086] = 6'b011101;
    assign data[2087] = 6'b011110;
    assign data[2088] = 6'b011110;
    assign data[2089] = 6'b011110;
    assign data[2090] = 6'b011111;
    assign data[2091] = 6'b011111;
    assign data[2092] = 6'b100000;
    assign data[2093] = 6'b100000;
    assign data[2094] = 6'b100001;
    assign data[2095] = 6'b100001;
    assign data[2096] = 6'b100010;
    assign data[2097] = 6'b100010;
    assign data[2098] = 6'b100011;
    assign data[2099] = 6'b100011;
    assign data[2100] = 6'b100100;
    assign data[2101] = 6'b100101;
    assign data[2102] = 6'b100101;
    assign data[2103] = 6'b100110;
    assign data[2104] = 6'b100111;
    assign data[2105] = 6'b100111;
    assign data[2106] = 6'b101000;
    assign data[2107] = 6'b101001;
    assign data[2108] = 6'b101001;
    assign data[2109] = 6'b101010;
    assign data[2110] = 6'b101011;
    assign data[2111] = 6'b101100;
    assign data[2112] = 6'b101100;
    assign data[2113] = 6'b101101;
    assign data[2114] = 6'b101110;
    assign data[2115] = 6'b011011;
    assign data[2116] = 6'b011011;
    assign data[2117] = 6'b011011;
    assign data[2118] = 6'b011100;
    assign data[2119] = 6'b011100;
    assign data[2120] = 6'b011100;
    assign data[2121] = 6'b011100;
    assign data[2122] = 6'b011100;
    assign data[2123] = 6'b011100;
    assign data[2124] = 6'b011100;
    assign data[2125] = 6'b011101;
    assign data[2126] = 6'b011101;
    assign data[2127] = 6'b011101;
    assign data[2128] = 6'b011101;
    assign data[2129] = 6'b011110;
    assign data[2130] = 6'b011110;
    assign data[2131] = 6'b011110;
    assign data[2132] = 6'b011111;
    assign data[2133] = 6'b011111;
    assign data[2134] = 6'b011111;
    assign data[2135] = 6'b100000;
    assign data[2136] = 6'b100000;
    assign data[2137] = 6'b100001;
    assign data[2138] = 6'b100001;
    assign data[2139] = 6'b100010;
    assign data[2140] = 6'b100010;
    assign data[2141] = 6'b100011;
    assign data[2142] = 6'b100011;
    assign data[2143] = 6'b100100;
    assign data[2144] = 6'b100100;
    assign data[2145] = 6'b100101;
    assign data[2146] = 6'b100101;
    assign data[2147] = 6'b100110;
    assign data[2148] = 6'b100111;
    assign data[2149] = 6'b100111;
    assign data[2150] = 6'b101000;
    assign data[2151] = 6'b101001;
    assign data[2152] = 6'b101001;
    assign data[2153] = 6'b101010;
    assign data[2154] = 6'b101011;
    assign data[2155] = 6'b101100;
    assign data[2156] = 6'b101100;
    assign data[2157] = 6'b101101;
    assign data[2158] = 6'b101110;
    assign data[2159] = 6'b101111;
    assign data[2160] = 6'b011100;
    assign data[2161] = 6'b011100;
    assign data[2162] = 6'b011101;
    assign data[2163] = 6'b011101;
    assign data[2164] = 6'b011101;
    assign data[2165] = 6'b011101;
    assign data[2166] = 6'b011101;
    assign data[2167] = 6'b011101;
    assign data[2168] = 6'b011101;
    assign data[2169] = 6'b011101;
    assign data[2170] = 6'b011110;
    assign data[2171] = 6'b011110;
    assign data[2172] = 6'b011110;
    assign data[2173] = 6'b011110;
    assign data[2174] = 6'b011111;
    assign data[2175] = 6'b011111;
    assign data[2176] = 6'b011111;
    assign data[2177] = 6'b100000;
    assign data[2178] = 6'b100000;
    assign data[2179] = 6'b100000;
    assign data[2180] = 6'b100001;
    assign data[2181] = 6'b100001;
    assign data[2182] = 6'b100010;
    assign data[2183] = 6'b100010;
    assign data[2184] = 6'b100011;
    assign data[2185] = 6'b100011;
    assign data[2186] = 6'b100100;
    assign data[2187] = 6'b100100;
    assign data[2188] = 6'b100101;
    assign data[2189] = 6'b100101;
    assign data[2190] = 6'b100110;
    assign data[2191] = 6'b100110;
    assign data[2192] = 6'b100111;
    assign data[2193] = 6'b101000;
    assign data[2194] = 6'b101000;
    assign data[2195] = 6'b101001;
    assign data[2196] = 6'b101010;
    assign data[2197] = 6'b101010;
    assign data[2198] = 6'b101011;
    assign data[2199] = 6'b101100;
    assign data[2200] = 6'b101100;
    assign data[2201] = 6'b101101;
    assign data[2202] = 6'b101110;
    assign data[2203] = 6'b101111;
    assign data[2204] = 6'b110000;
    assign data[2205] = 6'b011101;
    assign data[2206] = 6'b011101;
    assign data[2207] = 6'b011110;
    assign data[2208] = 6'b011110;
    assign data[2209] = 6'b011110;
    assign data[2210] = 6'b011110;
    assign data[2211] = 6'b011110;
    assign data[2212] = 6'b011110;
    assign data[2213] = 6'b011110;
    assign data[2214] = 6'b011110;
    assign data[2215] = 6'b011111;
    assign data[2216] = 6'b011111;
    assign data[2217] = 6'b011111;
    assign data[2218] = 6'b011111;
    assign data[2219] = 6'b100000;
    assign data[2220] = 6'b100000;
    assign data[2221] = 6'b100000;
    assign data[2222] = 6'b100001;
    assign data[2223] = 6'b100001;
    assign data[2224] = 6'b100001;
    assign data[2225] = 6'b100010;
    assign data[2226] = 6'b100010;
    assign data[2227] = 6'b100011;
    assign data[2228] = 6'b100011;
    assign data[2229] = 6'b100100;
    assign data[2230] = 6'b100100;
    assign data[2231] = 6'b100101;
    assign data[2232] = 6'b100101;
    assign data[2233] = 6'b100110;
    assign data[2234] = 6'b100110;
    assign data[2235] = 6'b100111;
    assign data[2236] = 6'b100111;
    assign data[2237] = 6'b101000;
    assign data[2238] = 6'b101001;
    assign data[2239] = 6'b101001;
    assign data[2240] = 6'b101010;
    assign data[2241] = 6'b101011;
    assign data[2242] = 6'b101011;
    assign data[2243] = 6'b101100;
    assign data[2244] = 6'b101101;
    assign data[2245] = 6'b101101;
    assign data[2246] = 6'b101110;
    assign data[2247] = 6'b101111;
    assign data[2248] = 6'b110000;
    assign data[2249] = 6'b110000;
    assign data[2250] = 6'b011111;
    assign data[2251] = 6'b011111;
    assign data[2252] = 6'b011111;
    assign data[2253] = 6'b011111;
    assign data[2254] = 6'b011111;
    assign data[2255] = 6'b011111;
    assign data[2256] = 6'b011111;
    assign data[2257] = 6'b011111;
    assign data[2258] = 6'b011111;
    assign data[2259] = 6'b011111;
    assign data[2260] = 6'b100000;
    assign data[2261] = 6'b100000;
    assign data[2262] = 6'b100000;
    assign data[2263] = 6'b100000;
    assign data[2264] = 6'b100001;
    assign data[2265] = 6'b100001;
    assign data[2266] = 6'b100001;
    assign data[2267] = 6'b100010;
    assign data[2268] = 6'b100010;
    assign data[2269] = 6'b100010;
    assign data[2270] = 6'b100011;
    assign data[2271] = 6'b100011;
    assign data[2272] = 6'b100100;
    assign data[2273] = 6'b100100;
    assign data[2274] = 6'b100101;
    assign data[2275] = 6'b100101;
    assign data[2276] = 6'b100110;
    assign data[2277] = 6'b100110;
    assign data[2278] = 6'b100111;
    assign data[2279] = 6'b100111;
    assign data[2280] = 6'b101000;
    assign data[2281] = 6'b101000;
    assign data[2282] = 6'b101001;
    assign data[2283] = 6'b101010;
    assign data[2284] = 6'b101010;
    assign data[2285] = 6'b101011;
    assign data[2286] = 6'b101011;
    assign data[2287] = 6'b101100;
    assign data[2288] = 6'b101101;
    assign data[2289] = 6'b101110;
    assign data[2290] = 6'b101110;
    assign data[2291] = 6'b101111;
    assign data[2292] = 6'b110000;
    assign data[2293] = 6'b110001;
    assign data[2294] = 6'b110001;
    assign data[2295] = 6'b100000;
    assign data[2296] = 6'b100000;
    assign data[2297] = 6'b100000;
    assign data[2298] = 6'b100000;
    assign data[2299] = 6'b100000;
    assign data[2300] = 6'b100000;
    assign data[2301] = 6'b100000;
    assign data[2302] = 6'b100000;
    assign data[2303] = 6'b100000;
    assign data[2304] = 6'b100000;
    assign data[2305] = 6'b100001;
    assign data[2306] = 6'b100001;
    assign data[2307] = 6'b100001;
    assign data[2308] = 6'b100001;
    assign data[2309] = 6'b100010;
    assign data[2310] = 6'b100010;
    assign data[2311] = 6'b100010;
    assign data[2312] = 6'b100011;
    assign data[2313] = 6'b100011;
    assign data[2314] = 6'b100011;
    assign data[2315] = 6'b100100;
    assign data[2316] = 6'b100100;
    assign data[2317] = 6'b100101;
    assign data[2318] = 6'b100101;
    assign data[2319] = 6'b100110;
    assign data[2320] = 6'b100110;
    assign data[2321] = 6'b100111;
    assign data[2322] = 6'b100111;
    assign data[2323] = 6'b101000;
    assign data[2324] = 6'b101000;
    assign data[2325] = 6'b101001;
    assign data[2326] = 6'b101001;
    assign data[2327] = 6'b101010;
    assign data[2328] = 6'b101010;
    assign data[2329] = 6'b101011;
    assign data[2330] = 6'b101100;
    assign data[2331] = 6'b101100;
    assign data[2332] = 6'b101101;
    assign data[2333] = 6'b101110;
    assign data[2334] = 6'b101110;
    assign data[2335] = 6'b101111;
    assign data[2336] = 6'b110000;
    assign data[2337] = 6'b110001;
    assign data[2338] = 6'b110001;
    assign data[2339] = 6'b110010;
    assign data[2340] = 6'b100001;
    assign data[2341] = 6'b100001;
    assign data[2342] = 6'b100001;
    assign data[2343] = 6'b100001;
    assign data[2344] = 6'b100001;
    assign data[2345] = 6'b100001;
    assign data[2346] = 6'b100001;
    assign data[2347] = 6'b100001;
    assign data[2348] = 6'b100001;
    assign data[2349] = 6'b100010;
    assign data[2350] = 6'b100010;
    assign data[2351] = 6'b100010;
    assign data[2352] = 6'b100010;
    assign data[2353] = 6'b100010;
    assign data[2354] = 6'b100011;
    assign data[2355] = 6'b100011;
    assign data[2356] = 6'b100011;
    assign data[2357] = 6'b100100;
    assign data[2358] = 6'b100100;
    assign data[2359] = 6'b100100;
    assign data[2360] = 6'b100101;
    assign data[2361] = 6'b100101;
    assign data[2362] = 6'b100110;
    assign data[2363] = 6'b100110;
    assign data[2364] = 6'b100111;
    assign data[2365] = 6'b100111;
    assign data[2366] = 6'b101000;
    assign data[2367] = 6'b101000;
    assign data[2368] = 6'b101001;
    assign data[2369] = 6'b101001;
    assign data[2370] = 6'b101010;
    assign data[2371] = 6'b101010;
    assign data[2372] = 6'b101011;
    assign data[2373] = 6'b101011;
    assign data[2374] = 6'b101100;
    assign data[2375] = 6'b101101;
    assign data[2376] = 6'b101101;
    assign data[2377] = 6'b101110;
    assign data[2378] = 6'b101111;
    assign data[2379] = 6'b101111;
    assign data[2380] = 6'b110000;
    assign data[2381] = 6'b110001;
    assign data[2382] = 6'b110010;
    assign data[2383] = 6'b110010;
    assign data[2384] = 6'b110011;
    assign data[2385] = 6'b100010;
    assign data[2386] = 6'b100010;
    assign data[2387] = 6'b100010;
    assign data[2388] = 6'b100010;
    assign data[2389] = 6'b100010;
    assign data[2390] = 6'b100010;
    assign data[2391] = 6'b100010;
    assign data[2392] = 6'b100010;
    assign data[2393] = 6'b100010;
    assign data[2394] = 6'b100011;
    assign data[2395] = 6'b100011;
    assign data[2396] = 6'b100011;
    assign data[2397] = 6'b100011;
    assign data[2398] = 6'b100100;
    assign data[2399] = 6'b100100;
    assign data[2400] = 6'b100100;
    assign data[2401] = 6'b100100;
    assign data[2402] = 6'b100101;
    assign data[2403] = 6'b100101;
    assign data[2404] = 6'b100101;
    assign data[2405] = 6'b100110;
    assign data[2406] = 6'b100110;
    assign data[2407] = 6'b100111;
    assign data[2408] = 6'b100111;
    assign data[2409] = 6'b101000;
    assign data[2410] = 6'b101000;
    assign data[2411] = 6'b101001;
    assign data[2412] = 6'b101001;
    assign data[2413] = 6'b101010;
    assign data[2414] = 6'b101010;
    assign data[2415] = 6'b101011;
    assign data[2416] = 6'b101011;
    assign data[2417] = 6'b101100;
    assign data[2418] = 6'b101100;
    assign data[2419] = 6'b101101;
    assign data[2420] = 6'b101110;
    assign data[2421] = 6'b101110;
    assign data[2422] = 6'b101111;
    assign data[2423] = 6'b110000;
    assign data[2424] = 6'b110000;
    assign data[2425] = 6'b110001;
    assign data[2426] = 6'b110010;
    assign data[2427] = 6'b110011;
    assign data[2428] = 6'b110011;
    assign data[2429] = 6'b110100;
    assign data[2430] = 6'b100011;
    assign data[2431] = 6'b100011;
    assign data[2432] = 6'b100011;
    assign data[2433] = 6'b100011;
    assign data[2434] = 6'b100011;
    assign data[2435] = 6'b100011;
    assign data[2436] = 6'b100011;
    assign data[2437] = 6'b100011;
    assign data[2438] = 6'b100011;
    assign data[2439] = 6'b100100;
    assign data[2440] = 6'b100100;
    assign data[2441] = 6'b100100;
    assign data[2442] = 6'b100100;
    assign data[2443] = 6'b100101;
    assign data[2444] = 6'b100101;
    assign data[2445] = 6'b100101;
    assign data[2446] = 6'b100101;
    assign data[2447] = 6'b100110;
    assign data[2448] = 6'b100110;
    assign data[2449] = 6'b100110;
    assign data[2450] = 6'b100111;
    assign data[2451] = 6'b100111;
    assign data[2452] = 6'b101000;
    assign data[2453] = 6'b101000;
    assign data[2454] = 6'b101001;
    assign data[2455] = 6'b101001;
    assign data[2456] = 6'b101010;
    assign data[2457] = 6'b101010;
    assign data[2458] = 6'b101011;
    assign data[2459] = 6'b101011;
    assign data[2460] = 6'b101100;
    assign data[2461] = 6'b101100;
    assign data[2462] = 6'b101101;
    assign data[2463] = 6'b101101;
    assign data[2464] = 6'b101110;
    assign data[2465] = 6'b101111;
    assign data[2466] = 6'b101111;
    assign data[2467] = 6'b110000;
    assign data[2468] = 6'b110001;
    assign data[2469] = 6'b110001;
    assign data[2470] = 6'b110010;
    assign data[2471] = 6'b110011;
    assign data[2472] = 6'b110011;
    assign data[2473] = 6'b110100;
    assign data[2474] = 6'b110101;

    Coordinate_generator c0(
        .p_x(p_x),
        .p_y(p_y),
        .real_x(real_x),
        .real_y(real_y)
    );

    genvar idx;
    generate
        for(idx=0; idx<16; idx=idx+1) begin: genXY
            abs_X x0(
                .x(real_x[idx]),
                .abs_real_x(abs_real_x[idx])
            );
            abs_Y y0(
                .y(real_y[idx]),
                .abs_real_y(abs_real_y[idx])
            );
            assign delta[idx] = `DELTA_START + data[abs_real_x[idx]*45+abs_real_y[idx]];
        end
    endgenerate



endmodule